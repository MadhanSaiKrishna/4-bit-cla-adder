magic
tech scmos
timestamp 1732037783
<< nwell >>
rect -420 33 -379 132
rect -340 33 -315 132
rect -281 34 -256 133
rect -225 78 -201 130
<< ntransistor >>
rect -214 47 -212 67
rect -408 -29 -406 11
rect -328 -29 -326 11
rect -269 -28 -267 12
rect -328 -103 -326 -63
rect -269 -102 -267 -62
<< ptransistor >>
rect -408 41 -406 121
rect -392 41 -390 121
rect -328 41 -326 121
rect -269 42 -267 122
rect -214 84 -212 124
<< ndiffusion >>
rect -215 47 -214 67
rect -212 47 -211 67
rect -409 -29 -408 11
rect -406 -29 -405 11
rect -329 -29 -328 11
rect -326 -29 -325 11
rect -270 -28 -269 12
rect -267 -28 -266 12
rect -329 -103 -328 -63
rect -326 -103 -325 -63
rect -270 -102 -269 -62
rect -267 -102 -266 -62
<< pdiffusion >>
rect -409 41 -408 121
rect -406 41 -405 121
rect -393 41 -392 121
rect -390 41 -389 121
rect -329 41 -328 121
rect -326 41 -325 121
rect -270 42 -269 122
rect -267 42 -266 122
rect -215 84 -214 124
rect -212 84 -211 124
<< ndcontact >>
rect -219 47 -215 67
rect -211 47 -207 67
rect -413 -29 -409 11
rect -405 -29 -401 11
rect -333 -29 -329 11
rect -325 -29 -321 11
rect -274 -28 -270 12
rect -266 -28 -262 12
rect -333 -103 -329 -63
rect -325 -103 -321 -63
rect -274 -102 -270 -62
rect -266 -102 -262 -62
<< pdcontact >>
rect -413 41 -409 121
rect -405 41 -401 121
rect -397 41 -393 121
rect -389 41 -385 121
rect -333 41 -329 121
rect -325 41 -321 121
rect -274 42 -270 122
rect -266 42 -262 122
rect -219 84 -215 124
rect -211 84 -207 124
<< polysilicon >>
rect -408 121 -406 125
rect -392 121 -390 125
rect -328 121 -326 125
rect -269 122 -267 126
rect -214 124 -212 130
rect -214 67 -212 84
rect -214 43 -212 47
rect -408 11 -406 41
rect -392 19 -390 41
rect -328 32 -326 41
rect -269 29 -267 42
rect -328 11 -326 14
rect -269 12 -267 15
rect -408 -33 -406 -29
rect -328 -33 -326 -29
rect -269 -35 -267 -28
rect -328 -63 -326 -56
rect -269 -62 -267 -55
rect -328 -107 -326 -103
rect -269 -106 -267 -102
<< polycontact >>
rect -219 71 -214 75
rect -414 23 -408 28
rect -390 22 -385 27
rect -329 22 -325 32
rect -271 22 -264 29
rect -329 14 -325 18
rect -271 -40 -264 -35
rect -331 -56 -326 -51
rect -272 -55 -267 -50
<< metal1 >>
rect -420 129 -315 135
rect -413 121 -409 129
rect -340 127 -315 129
rect -281 128 -256 136
rect -225 130 -201 134
rect -333 121 -329 127
rect -274 122 -270 128
rect -219 124 -215 130
rect -401 41 -397 121
rect -385 47 -381 121
rect -385 41 -373 47
rect -380 34 -373 41
rect -380 31 -346 34
rect -391 22 -390 27
rect -380 11 -373 31
rect -349 18 -346 31
rect -321 29 -315 121
rect -262 89 -256 122
rect -262 84 -242 89
rect -262 42 -256 84
rect -247 75 -242 84
rect -211 75 -207 84
rect -247 71 -219 75
rect -211 71 -201 75
rect -321 22 -271 29
rect -264 22 -263 29
rect -349 14 -329 18
rect -401 5 -373 11
rect -401 -29 -400 5
rect -321 -3 -315 22
rect -288 -2 -274 4
rect -413 -33 -409 -29
rect -423 -40 -379 -33
rect -333 -51 -329 -29
rect -333 -56 -331 -51
rect -333 -63 -329 -56
rect -288 -77 -284 -2
rect -247 4 -242 71
rect -211 67 -207 71
rect -219 43 -214 47
rect -225 39 -201 43
rect -262 -2 -242 4
rect -274 -32 -270 -28
rect -288 -84 -274 -77
rect -325 -107 -321 -103
rect -266 -106 -262 -102
rect -338 -113 -310 -107
rect -279 -112 -251 -106
<< m2contact >>
rect -263 22 -256 29
<< metal2 >>
rect -419 23 -408 28
rect -391 22 -325 27
rect -256 22 -228 29
rect -358 -35 -355 22
rect -358 -40 -264 -35
rect -358 -51 -355 -40
rect -235 -50 -228 22
rect -358 -56 -326 -51
rect -267 -55 -228 -50
<< labels >>
rlabel metal1 -270 133 -270 133 5 vdd
rlabel metal1 -266 -108 -266 -108 1 gnd
rlabel metal2 -384 24 -384 24 1 clk
rlabel metal1 -376 33 -376 33 1 n1
rlabel metal1 -329 132 -329 132 5 vdd
rlabel metal1 -325 -109 -325 -109 1 gnd
rlabel metal2 -417 26 -417 26 1 a_in
rlabel metal1 -405 -37 -405 -37 1 gnd
rlabel metal1 -400 133 -400 133 5 vdd
rlabel metal1 -214 41 -214 41 1 gnd
rlabel metal1 -214 132 -214 132 5 vdd
rlabel metal1 -242 73 -242 73 1 n3
rlabel metal1 -207 72 -205 74 7 a
rlabel metal1 -222 73 -222 73 3 in
rlabel metal1 -310 25 -310 25 1 n2
<< end >>
