magic
tech scmos
timestamp 1733164831
<< nwell >>
rect 21 97 45 149
rect 65 57 125 149
rect -18 -10 6 42
<< ntransistor >>
rect 32 66 34 86
rect -7 -41 -5 -21
rect 76 -42 78 -2
rect 88 -42 90 -2
rect 100 -42 102 -2
rect 112 -42 114 -2
<< ptransistor >>
rect 32 103 34 143
rect 76 63 78 143
rect 88 63 90 143
rect 100 63 102 143
rect 112 63 114 143
rect -7 -4 -5 36
<< ndiffusion >>
rect 31 66 32 86
rect 34 66 35 86
rect -8 -41 -7 -21
rect -5 -41 -4 -21
rect 75 -42 76 -2
rect 78 -42 79 -2
rect 87 -42 88 -2
rect 90 -42 91 -2
rect 99 -42 100 -2
rect 102 -40 103 -2
rect 111 -40 112 -2
rect 102 -42 112 -40
rect 114 -42 115 -2
<< pdiffusion >>
rect 31 103 32 143
rect 34 103 35 143
rect 75 63 76 143
rect 78 63 79 143
rect 87 63 88 143
rect 90 63 91 143
rect 99 63 100 143
rect 102 63 103 143
rect 111 63 112 143
rect 114 63 115 143
rect -8 -4 -7 36
rect -5 -4 -4 36
<< ndcontact >>
rect 27 66 31 86
rect 35 66 39 86
rect -12 -41 -8 -21
rect -4 -41 0 -21
rect 71 -42 75 -2
rect 79 -42 87 -2
rect 91 -42 99 -2
rect 103 -40 111 -2
rect 115 -42 119 -2
<< pdcontact >>
rect 27 103 31 143
rect 35 103 39 143
rect 71 63 75 143
rect 79 63 87 143
rect 91 63 99 143
rect 103 63 111 143
rect 115 63 119 143
rect -12 -4 -8 36
rect -4 -4 0 36
<< polysilicon >>
rect 32 143 34 149
rect 76 143 78 147
rect 88 143 90 147
rect 100 143 102 147
rect 112 143 114 147
rect 32 86 34 103
rect 32 62 34 66
rect -7 36 -5 42
rect 76 -2 78 63
rect 88 -2 90 63
rect 100 -2 102 63
rect 112 -2 114 63
rect -7 -21 -5 -4
rect -7 -45 -5 -41
rect 76 -46 78 -42
rect 88 -46 90 -42
rect 100 -47 102 -42
rect 112 -47 114 -42
<< polycontact >>
rect 27 90 32 94
rect 70 40 76 44
rect 83 32 88 36
rect 95 22 100 26
rect 108 12 112 16
rect -12 -17 -7 -13
<< metal1 >>
rect -12 149 125 153
rect -30 90 -20 94
rect -12 36 -8 149
rect 27 143 31 149
rect 91 143 99 149
rect 35 94 39 103
rect 6 90 27 94
rect 35 90 50 94
rect 7 28 12 90
rect 35 86 39 90
rect -28 -17 -24 -13
rect -4 -13 0 -4
rect -19 -17 -12 -13
rect -4 -17 15 -13
rect -4 -21 0 -17
rect -12 -49 -8 -41
rect 27 -49 31 66
rect 46 44 50 90
rect 71 55 75 63
rect 115 55 119 63
rect 71 50 135 55
rect 46 40 70 44
rect 54 32 83 36
rect 53 22 95 26
rect 46 12 108 16
rect 46 -12 51 12
rect 71 2 119 7
rect 71 -2 75 2
rect 115 -2 119 2
rect 103 -42 111 -40
rect 81 -49 85 -42
rect -12 -53 85 -49
rect 105 -49 109 -42
rect 123 -49 127 50
rect 105 -53 127 -49
<< m2contact >>
rect -20 89 -15 95
rect 1 90 6 95
rect 7 21 13 28
rect -24 -17 -19 -12
rect 15 -18 21 -12
rect 48 31 54 37
rect 47 20 53 27
rect 45 -17 51 -12
<< metal2 >>
rect -15 90 1 94
rect -23 32 48 36
rect -23 -12 -19 32
rect 13 22 47 26
rect 21 -17 45 -13
<< labels >>
rlabel metal1 132 53 132 53 1 P0
rlabel metal1 -7 -51 -7 -51 1 gnd
rlabel metal1 -7 151 -7 151 5 vdd
rlabel metal1 34 -51 34 -51 1 gnd
rlabel metal1 32 152 32 152 5 vdd
rlabel space -18 -18 -12 -13 1 a0
rlabel space -2 -18 5 -11 1 a0_inv
rlabel metal1 40 90 46 94 1 b0_inv
rlabel metal1 103 13 107 16 1 a0_inv
rlabel metal1 91 23 95 26 1 b0
rlabel metal1 78 32 82 35 1 a0
rlabel metal1 65 41 69 44 1 b0_inv
rlabel metal1 15 90 22 94 1 b0
rlabel space -27 90 -20 96 1 b0
<< end >>
