.include inverter.cir
.subckt cpl_dff b_in b clk vdd gnd

.param width_P = 40*LAMBDA
.param width_N = 20*LAMBDA

M1 b_in clk n1 n1 CMOSN W={width_N} L={2*LAMBDA}
+AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+AD={5*width_N*LAMBDA} PD = {10*LAMBDA+2*width_N}

M2 n1 clk b_in b_in CMOSP W={width_P} L={2*LAMBDA}
+AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

X1 n1 n2 vdd gnd inverter width_P={width_P} width_N={width_N}
X2 n2 n1 vdd gnd inverter width_P ={width_P} width_N={width_N}

M3 n2 clk n3 n3 CMOSN W={width_N} L={2*LAMBDA}
+AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+AD={5*width_N*LAMBDA} PD = {10*LAMBDA+2*width_N}

M4 n3 clk n2 n2  CMOSP W={width_P} L={2*LAMBDA}
+AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

X3 n3 b vdd gnd inverter width_P={width_P} width_N={width_N}
X4 b n3 vdd gnd inverter width_P={width_P} width_N={width_N}

.ends cpl_dff