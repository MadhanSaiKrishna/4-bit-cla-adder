magic
tech scmos
timestamp 1733176363
<< nwell >>
rect 349 81 458 214
rect 471 81 496 214
rect 568 53 592 105
<< ntransistor >>
rect 579 22 581 42
rect 360 -117 362 -57
rect 372 -117 374 -57
rect 384 -117 386 -57
rect 396 -117 398 -57
rect 408 -117 410 -57
rect 420 -117 422 -57
rect 432 -117 434 -57
rect 444 -117 446 -57
rect 482 -118 484 -57
<< ptransistor >>
rect 360 87 362 207
rect 372 87 374 207
rect 384 87 386 207
rect 396 87 398 207
rect 408 87 410 207
rect 420 87 422 207
rect 432 87 434 207
rect 444 87 446 207
rect 482 87 484 207
rect 579 59 581 99
<< ndiffusion >>
rect 578 22 579 42
rect 581 22 582 42
rect 359 -117 360 -57
rect 362 -117 363 -57
rect 371 -117 372 -57
rect 374 -117 375 -57
rect 383 -117 384 -57
rect 386 -117 387 -57
rect 395 -117 396 -57
rect 398 -117 399 -57
rect 407 -117 408 -57
rect 410 -117 411 -57
rect 419 -117 420 -57
rect 422 -117 423 -57
rect 431 -117 432 -57
rect 434 -117 435 -57
rect 443 -117 444 -57
rect 446 -117 447 -57
rect 481 -118 482 -57
rect 484 -118 485 -57
<< pdiffusion >>
rect 359 87 360 207
rect 362 87 363 207
rect 371 87 372 207
rect 374 87 375 207
rect 383 87 384 207
rect 386 87 387 207
rect 395 87 396 207
rect 398 87 399 207
rect 407 87 408 207
rect 410 87 411 207
rect 419 87 420 207
rect 422 87 423 207
rect 431 87 432 207
rect 434 87 435 207
rect 443 87 444 207
rect 446 87 447 207
rect 481 87 482 207
rect 484 87 485 207
rect 578 59 579 99
rect 581 59 582 99
<< ndcontact >>
rect 574 22 578 42
rect 582 22 586 42
rect 355 -117 359 -57
rect 363 -117 371 -57
rect 375 -117 383 -57
rect 387 -117 395 -57
rect 399 -117 407 -57
rect 411 -117 419 -57
rect 423 -117 431 -57
rect 435 -117 443 -57
rect 447 -117 451 -57
rect 477 -118 481 -57
rect 485 -118 489 -57
<< pdcontact >>
rect 355 87 359 207
rect 363 87 371 207
rect 375 87 383 207
rect 387 87 395 207
rect 399 87 407 207
rect 411 87 419 207
rect 423 87 431 207
rect 435 87 443 207
rect 447 87 451 207
rect 477 87 481 207
rect 485 87 489 207
rect 574 59 578 99
rect 582 59 586 99
<< polysilicon >>
rect 360 207 362 210
rect 372 207 374 210
rect 384 207 386 210
rect 396 207 398 210
rect 408 207 410 210
rect 420 207 422 210
rect 432 207 434 210
rect 444 207 446 210
rect 482 207 484 210
rect 579 99 581 105
rect 360 23 362 87
rect 372 23 374 87
rect 360 -57 362 19
rect 372 -57 374 19
rect 384 -57 386 87
rect 396 -57 398 87
rect 408 -57 410 87
rect 420 -57 422 87
rect 432 -57 434 87
rect 444 -57 446 87
rect 482 -57 484 87
rect 579 42 581 59
rect 579 18 581 22
rect 360 -125 362 -117
rect 372 -125 374 -117
rect 384 -126 386 -117
rect 396 -126 398 -117
rect 408 -126 410 -117
rect 420 -125 422 -117
rect 432 -125 434 -117
rect 444 -125 446 -117
rect 482 -125 484 -118
<< polycontact >>
rect 356 36 360 40
rect 368 27 372 31
rect 380 19 384 23
rect 392 11 396 15
rect 404 3 408 7
rect 416 -5 420 -1
rect 428 -15 432 -11
rect 440 -23 444 -19
rect 478 -31 482 -27
rect 574 46 579 50
<< metal1 >>
rect 355 223 577 227
rect 355 207 359 223
rect 413 207 417 223
rect 425 215 481 218
rect 425 207 429 215
rect 477 207 481 215
rect 377 51 380 87
rect 389 58 392 87
rect 438 58 441 87
rect 447 76 450 87
rect 485 58 489 87
rect 574 99 577 223
rect 389 55 489 58
rect 381 47 447 50
rect 582 50 586 59
rect 452 47 574 50
rect 582 46 602 50
rect 377 44 380 46
rect 582 42 586 46
rect 326 36 336 40
rect 342 36 356 40
rect 326 27 368 31
rect 355 23 358 27
rect 355 19 380 23
rect 327 11 364 15
rect 369 11 392 15
rect 327 3 347 7
rect 352 3 404 7
rect 327 -5 416 -1
rect 352 -15 428 -11
rect 342 -23 440 -19
rect 369 -31 478 -27
rect 389 -41 489 -38
rect 377 -57 380 -42
rect 389 -57 392 -41
rect 437 -57 440 -41
rect 447 -57 450 -49
rect 486 -57 489 -41
rect 355 -135 359 -117
rect 426 -127 429 -117
rect 477 -127 480 -118
rect 426 -130 480 -127
rect 574 -135 578 22
rect 355 -140 578 -135
<< m2contact >>
rect 447 70 452 76
rect 376 46 381 51
rect 447 46 452 51
rect 336 36 342 41
rect 364 11 369 16
rect 347 3 352 8
rect 347 -15 352 -10
rect 336 -23 342 -18
rect 364 -31 369 -26
rect 376 -42 381 -37
rect 447 -49 452 -44
<< metal2 >>
rect 447 51 450 70
rect 337 -18 342 36
rect 377 23 380 46
rect 348 -10 352 3
rect 365 -26 369 11
rect 377 -37 380 19
rect 447 -44 450 46
rect 447 -57 450 -49
<< labels >>
rlabel metal1 384 224 388 226 5 vdd
rlabel metal1 567 224 576 227 5 vdd
rlabel metal1 382 -139 388 -137 1 gnd
rlabel metal1 328 27 334 31 3 b1
rlabel metal1 326 36 333 40 3 a1
rlabel metal1 330 11 336 15 1 b0
rlabel metal1 331 -5 336 -1 1 cin
rlabel metal1 330 3 335 7 1 a0
rlabel metal1 566 -139 573 -136 1 gnd
rlabel metal1 590 46 595 50 1 c2
<< end >>
