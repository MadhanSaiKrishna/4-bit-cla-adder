.subckt two_xor a0 b0 p0 vdd gnd

.param width_P = 40*LAMBDA
.param width_N = 20*LAMBDA

M1 a0_inv a0 vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M2 a0_inv a0 gnd gnd CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M3 b0_inv b0 vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M4 b0_inv b0 gnd gnd CMOSN W={width_N} L={2*LAMBDA} 
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M5 n1 a0 vdd vdd CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

M6 p0 b0_inv n1 n1 CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

M7 p0 b0 n2 n2 CMOSN W={2*width_N} L={2*LAMBDA} 
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N}
+ AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*2*width_N}

M8 n2 a0 gnd gnd CMOSN W={2*width_N} L={2*LAMBDA} 
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N}
+ AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*2*width_N}

M9 n3 b0 vdd vdd CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

M10 p0 a0_inv n3 n3 CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

M11 p0 b0_inv n4 n4 CMOSN W={2*width_N} L={2*LAMBDA} 
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N}
+ AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*2*width_N}

M12 n4 a0_inv gnd gnd CMOSN W={2*width_N} L={2*LAMBDA} 
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N}
+ AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*2*width_N}

.ends