magic
tech scmos
timestamp 1733242492
<< nwell >>
rect 692 883 889 936
rect 902 883 927 936
rect 941 883 966 936
rect 985 824 1009 876
rect 1297 648 1321 700
rect 1341 608 1401 700
rect 1469 648 1493 700
rect 1513 608 1573 700
rect 1258 541 1282 593
rect 1430 541 1454 593
rect 686 449 831 502
rect 844 449 869 502
rect 883 449 908 502
rect 919 379 943 431
rect 1292 360 1316 412
rect 1336 320 1396 412
rect 1464 360 1488 412
rect 1508 320 1568 412
rect 1253 253 1277 305
rect 1425 253 1449 305
rect -189 88 -152 187
rect -139 90 -113 187
rect -93 90 -67 187
rect -61 91 -33 143
rect -21 88 16 187
rect 29 90 55 187
rect 75 90 101 187
rect 107 91 135 143
rect 145 88 182 187
rect 195 90 221 187
rect 241 90 267 187
rect 273 91 301 143
rect 310 88 347 187
rect 360 90 386 187
rect 406 90 432 187
rect 438 91 466 143
rect 687 31 795 83
rect 812 31 836 83
rect 1290 71 1314 123
rect 868 14 892 66
rect 1334 31 1394 123
rect 1462 71 1486 123
rect 1506 31 1566 123
rect 1251 -36 1275 16
rect 1423 -36 1447 16
rect -190 -163 -153 -64
rect -140 -161 -114 -64
rect -94 -161 -68 -64
rect -62 -160 -34 -108
rect -22 -163 15 -64
rect 28 -161 54 -64
rect 74 -161 100 -64
rect 106 -160 134 -108
rect 144 -163 181 -64
rect 194 -161 220 -64
rect 240 -161 266 -64
rect 272 -160 300 -108
rect 309 -163 346 -64
rect 359 -161 385 -64
rect 405 -161 431 -64
rect 437 -160 465 -108
rect 1287 -236 1311 -184
rect 677 -314 743 -261
rect 749 -314 775 -261
rect 782 -313 806 -261
rect 1331 -276 1391 -184
rect 1459 -236 1483 -184
rect 1503 -276 1563 -184
rect 1248 -343 1272 -291
rect 1420 -343 1444 -291
<< ntransistor >>
rect 996 793 998 813
rect 1308 617 1310 637
rect 1480 617 1482 637
rect 707 551 709 571
rect 719 551 721 571
rect 731 551 733 571
rect 743 551 745 571
rect 755 551 757 571
rect 767 551 769 571
rect 779 551 781 571
rect 791 551 793 571
rect 803 551 805 571
rect 815 551 817 571
rect 827 551 829 571
rect 839 551 841 571
rect 851 551 853 571
rect 863 551 865 571
rect 875 551 877 571
rect 913 551 915 571
rect 952 551 954 571
rect 1269 510 1271 530
rect 1352 509 1354 549
rect 1364 509 1366 549
rect 1376 509 1378 549
rect 1388 509 1390 549
rect 1441 510 1443 530
rect 1524 509 1526 549
rect 1536 509 1538 549
rect 1548 509 1550 549
rect 1560 509 1562 549
rect 930 348 932 368
rect 1303 329 1305 349
rect 1475 329 1477 349
rect 1264 222 1266 242
rect 1347 221 1349 261
rect 1359 221 1361 261
rect 1371 221 1373 261
rect 1383 221 1385 261
rect 1436 222 1438 242
rect 1519 221 1521 261
rect 1531 221 1533 261
rect 1543 221 1545 261
rect 1555 221 1557 261
rect -46 60 -44 80
rect -177 12 -175 52
rect -126 15 -124 55
rect -114 15 -112 55
rect -80 15 -78 55
rect -68 15 -66 55
rect 122 60 124 80
rect -9 12 -7 52
rect 42 15 44 55
rect 54 15 56 55
rect 88 15 90 55
rect 100 15 102 55
rect 697 164 699 184
rect 709 164 711 184
rect 721 164 723 184
rect 733 164 735 184
rect 745 164 747 184
rect 757 164 759 184
rect 769 164 771 184
rect 781 164 783 184
rect 793 164 795 184
rect 805 164 807 184
rect 817 164 819 184
rect 855 164 857 184
rect 894 164 896 184
rect 288 60 290 80
rect 157 12 159 52
rect 208 15 210 55
rect 220 15 222 55
rect 254 15 256 55
rect 266 15 268 55
rect 453 60 455 80
rect 322 12 324 52
rect 373 15 375 55
rect 385 15 387 55
rect 419 15 421 55
rect 431 15 433 55
rect -47 -191 -45 -171
rect -178 -239 -176 -199
rect -127 -236 -125 -196
rect -115 -236 -113 -196
rect -81 -236 -79 -196
rect -69 -236 -67 -196
rect 121 -191 123 -171
rect -10 -239 -8 -199
rect 41 -236 43 -196
rect 53 -236 55 -196
rect 87 -236 89 -196
rect 99 -236 101 -196
rect 1301 40 1303 60
rect 1473 40 1475 60
rect 879 -17 881 3
rect 1262 -67 1264 -47
rect 1345 -68 1347 -28
rect 1357 -68 1359 -28
rect 1369 -68 1371 -28
rect 1381 -68 1383 -28
rect 1434 -67 1436 -47
rect 1517 -68 1519 -28
rect 1529 -68 1531 -28
rect 1541 -68 1543 -28
rect 1553 -68 1555 -28
rect 698 -101 700 -81
rect 710 -101 712 -81
rect 722 -101 724 -81
rect 734 -101 736 -81
rect 746 -101 748 -81
rect 758 -101 760 -81
rect 770 -101 772 -81
rect 782 -101 784 -81
rect 823 -101 825 -81
rect 287 -191 289 -171
rect 156 -239 158 -199
rect 207 -236 209 -196
rect 219 -236 221 -196
rect 253 -236 255 -196
rect 265 -236 267 -196
rect 452 -191 454 -171
rect 321 -239 323 -199
rect 372 -236 374 -196
rect 384 -236 386 -196
rect 418 -236 420 -196
rect 430 -236 432 -196
rect 1298 -267 1300 -247
rect 1470 -267 1472 -247
rect 688 -370 690 -350
rect 700 -370 702 -350
rect 712 -370 714 -350
rect 724 -370 726 -350
rect 761 -370 763 -350
rect 793 -393 795 -373
rect 1259 -374 1261 -354
rect 1342 -375 1344 -335
rect 1354 -375 1356 -335
rect 1366 -375 1368 -335
rect 1378 -375 1380 -335
rect 1431 -374 1433 -354
rect 1514 -375 1516 -335
rect 1526 -375 1528 -335
rect 1538 -375 1540 -335
rect 1550 -375 1552 -335
<< ptransistor >>
rect 707 889 709 929
rect 719 889 721 929
rect 731 889 733 929
rect 743 889 745 929
rect 755 889 757 929
rect 767 889 769 929
rect 779 889 781 929
rect 791 889 793 929
rect 803 889 805 929
rect 815 889 817 929
rect 827 889 829 929
rect 839 889 841 929
rect 851 889 853 929
rect 863 889 865 929
rect 875 889 877 929
rect 913 889 915 929
rect 952 889 954 929
rect 996 830 998 870
rect 1308 654 1310 694
rect 1352 614 1354 694
rect 1364 614 1366 694
rect 1376 614 1378 694
rect 1388 614 1390 694
rect 1480 654 1482 694
rect 1269 547 1271 587
rect 1524 614 1526 694
rect 1536 614 1538 694
rect 1548 614 1550 694
rect 1560 614 1562 694
rect 1441 547 1443 587
rect 697 455 699 495
rect 709 455 711 495
rect 721 455 723 495
rect 733 455 735 495
rect 745 455 747 495
rect 757 455 759 495
rect 769 455 771 495
rect 781 455 783 495
rect 793 455 795 495
rect 805 455 807 495
rect 817 455 819 495
rect 855 455 857 495
rect 894 455 896 495
rect 930 385 932 425
rect 1303 366 1305 406
rect 1347 326 1349 406
rect 1359 326 1361 406
rect 1371 326 1373 406
rect 1383 326 1385 406
rect 1475 366 1477 406
rect 1264 259 1266 299
rect 1519 326 1521 406
rect 1531 326 1533 406
rect 1543 326 1545 406
rect 1555 326 1557 406
rect 1436 259 1438 299
rect -177 96 -175 176
rect -165 96 -163 176
rect -126 96 -124 176
rect -80 96 -78 176
rect -46 97 -44 137
rect -9 96 -7 176
rect 3 96 5 176
rect 42 96 44 176
rect 88 96 90 176
rect 122 97 124 137
rect 157 96 159 176
rect 169 96 171 176
rect 208 96 210 176
rect 254 96 256 176
rect 288 97 290 137
rect 322 96 324 176
rect 334 96 336 176
rect 373 96 375 176
rect 419 96 421 176
rect 453 97 455 137
rect 1301 77 1303 117
rect 698 37 700 77
rect 710 37 712 77
rect 722 37 724 77
rect 734 37 736 77
rect 746 37 748 77
rect 758 37 760 77
rect 770 37 772 77
rect 782 37 784 77
rect 823 37 825 77
rect -178 -155 -176 -75
rect -166 -155 -164 -75
rect -127 -155 -125 -75
rect -81 -155 -79 -75
rect -47 -154 -45 -114
rect -10 -155 -8 -75
rect 2 -155 4 -75
rect 41 -155 43 -75
rect 87 -155 89 -75
rect 121 -154 123 -114
rect 156 -155 158 -75
rect 168 -155 170 -75
rect 207 -155 209 -75
rect 253 -155 255 -75
rect 287 -154 289 -114
rect 321 -155 323 -75
rect 333 -155 335 -75
rect 372 -155 374 -75
rect 418 -155 420 -75
rect 879 20 881 60
rect 1345 37 1347 117
rect 1357 37 1359 117
rect 1369 37 1371 117
rect 1381 37 1383 117
rect 1473 77 1475 117
rect 1262 -30 1264 10
rect 1517 37 1519 117
rect 1529 37 1531 117
rect 1541 37 1543 117
rect 1553 37 1555 117
rect 1434 -30 1436 10
rect 452 -154 454 -114
rect 1298 -230 1300 -190
rect 688 -308 690 -268
rect 700 -308 702 -268
rect 712 -308 714 -268
rect 724 -308 726 -268
rect 761 -308 763 -268
rect 793 -307 795 -267
rect 1342 -270 1344 -190
rect 1354 -270 1356 -190
rect 1366 -270 1368 -190
rect 1378 -270 1380 -190
rect 1470 -230 1472 -190
rect 1259 -337 1261 -297
rect 1514 -270 1516 -190
rect 1526 -270 1528 -190
rect 1538 -270 1540 -190
rect 1550 -270 1552 -190
rect 1431 -337 1433 -297
<< ndiffusion >>
rect 995 793 996 813
rect 998 793 999 813
rect 1307 617 1308 637
rect 1310 617 1311 637
rect 1479 617 1480 637
rect 1482 617 1483 637
rect 706 551 707 571
rect 709 551 710 571
rect 718 551 719 571
rect 721 551 722 571
rect 730 551 731 571
rect 733 551 734 571
rect 742 551 743 571
rect 745 551 746 571
rect 754 551 755 571
rect 757 551 758 571
rect 766 551 767 571
rect 769 551 770 571
rect 778 551 779 571
rect 781 551 782 571
rect 790 551 791 571
rect 793 551 794 571
rect 802 551 803 571
rect 805 551 806 571
rect 814 551 815 571
rect 817 551 818 571
rect 826 551 827 571
rect 829 551 830 571
rect 838 551 839 571
rect 841 551 842 571
rect 850 551 851 571
rect 853 551 854 571
rect 862 551 863 571
rect 865 551 866 571
rect 874 551 875 571
rect 877 551 878 571
rect 912 551 913 571
rect 915 551 916 571
rect 951 551 952 571
rect 954 551 955 571
rect 1268 510 1269 530
rect 1271 510 1272 530
rect 1351 509 1352 549
rect 1354 509 1355 549
rect 1363 509 1364 549
rect 1366 509 1367 549
rect 1375 509 1376 549
rect 1378 511 1379 549
rect 1387 511 1388 549
rect 1378 509 1388 511
rect 1390 509 1391 549
rect 1440 510 1441 530
rect 1443 510 1444 530
rect 1523 509 1524 549
rect 1526 509 1527 549
rect 1535 509 1536 549
rect 1538 509 1539 549
rect 1547 509 1548 549
rect 1550 511 1551 549
rect 1559 511 1560 549
rect 1550 509 1560 511
rect 1562 509 1563 549
rect 929 348 930 368
rect 932 348 933 368
rect 1302 329 1303 349
rect 1305 329 1306 349
rect 1474 329 1475 349
rect 1477 329 1478 349
rect 1263 222 1264 242
rect 1266 222 1267 242
rect 1346 221 1347 261
rect 1349 221 1350 261
rect 1358 221 1359 261
rect 1361 221 1362 261
rect 1370 221 1371 261
rect 1373 223 1374 261
rect 1382 223 1383 261
rect 1373 221 1383 223
rect 1385 221 1386 261
rect 1435 222 1436 242
rect 1438 222 1439 242
rect 1518 221 1519 261
rect 1521 221 1522 261
rect 1530 221 1531 261
rect 1533 221 1534 261
rect 1542 221 1543 261
rect 1545 223 1546 261
rect 1554 223 1555 261
rect 1545 221 1555 223
rect 1557 221 1558 261
rect -47 60 -46 80
rect -44 60 -43 80
rect -178 12 -177 52
rect -175 12 -174 52
rect -127 15 -126 55
rect -124 15 -123 55
rect -115 15 -114 55
rect -112 15 -111 55
rect -81 15 -80 55
rect -78 15 -77 55
rect -69 15 -68 55
rect -66 15 -65 55
rect 121 60 122 80
rect 124 60 125 80
rect -10 12 -9 52
rect -7 12 -6 52
rect 41 15 42 55
rect 44 15 45 55
rect 53 15 54 55
rect 56 15 57 55
rect 87 15 88 55
rect 90 15 91 55
rect 99 15 100 55
rect 102 15 103 55
rect 696 164 697 184
rect 699 164 700 184
rect 708 164 709 184
rect 711 164 712 184
rect 720 164 721 184
rect 723 164 724 184
rect 732 164 733 184
rect 735 164 736 184
rect 744 164 745 184
rect 747 164 748 184
rect 756 164 757 184
rect 759 164 760 184
rect 768 164 769 184
rect 771 164 772 184
rect 780 164 781 184
rect 783 164 784 184
rect 792 164 793 184
rect 795 164 796 184
rect 804 164 805 184
rect 807 164 808 184
rect 816 164 817 184
rect 819 164 820 184
rect 854 164 855 184
rect 857 164 858 184
rect 893 164 894 184
rect 896 164 897 184
rect 287 60 288 80
rect 290 60 291 80
rect 156 12 157 52
rect 159 12 160 52
rect 207 15 208 55
rect 210 15 211 55
rect 219 15 220 55
rect 222 15 223 55
rect 253 15 254 55
rect 256 15 257 55
rect 265 15 266 55
rect 268 15 269 55
rect 452 60 453 80
rect 455 60 456 80
rect 321 12 322 52
rect 324 12 325 52
rect 372 15 373 55
rect 375 15 376 55
rect 384 15 385 55
rect 387 15 388 55
rect 418 15 419 55
rect 421 15 422 55
rect 430 15 431 55
rect 433 15 434 55
rect -48 -191 -47 -171
rect -45 -191 -44 -171
rect -179 -239 -178 -199
rect -176 -239 -175 -199
rect -128 -236 -127 -196
rect -125 -236 -124 -196
rect -116 -236 -115 -196
rect -113 -236 -112 -196
rect -82 -236 -81 -196
rect -79 -236 -78 -196
rect -70 -236 -69 -196
rect -67 -236 -66 -196
rect 120 -191 121 -171
rect 123 -191 124 -171
rect -11 -239 -10 -199
rect -8 -239 -7 -199
rect 40 -236 41 -196
rect 43 -236 44 -196
rect 52 -236 53 -196
rect 55 -236 56 -196
rect 86 -236 87 -196
rect 89 -236 90 -196
rect 98 -236 99 -196
rect 101 -236 102 -196
rect 1300 40 1301 60
rect 1303 40 1304 60
rect 1472 40 1473 60
rect 1475 40 1476 60
rect 878 -17 879 3
rect 881 -17 882 3
rect 1261 -67 1262 -47
rect 1264 -67 1265 -47
rect 1344 -68 1345 -28
rect 1347 -68 1348 -28
rect 1356 -68 1357 -28
rect 1359 -68 1360 -28
rect 1368 -68 1369 -28
rect 1371 -66 1372 -28
rect 1380 -66 1381 -28
rect 1371 -68 1381 -66
rect 1383 -68 1384 -28
rect 1433 -67 1434 -47
rect 1436 -67 1437 -47
rect 1516 -68 1517 -28
rect 1519 -68 1520 -28
rect 1528 -68 1529 -28
rect 1531 -68 1532 -28
rect 1540 -68 1541 -28
rect 1543 -66 1544 -28
rect 1552 -66 1553 -28
rect 1543 -68 1553 -66
rect 1555 -68 1556 -28
rect 697 -101 698 -81
rect 700 -101 701 -81
rect 709 -101 710 -81
rect 712 -101 713 -81
rect 721 -101 722 -81
rect 724 -101 725 -81
rect 733 -101 734 -81
rect 736 -101 737 -81
rect 745 -101 746 -81
rect 748 -101 749 -81
rect 757 -101 758 -81
rect 760 -101 761 -81
rect 769 -101 770 -81
rect 772 -101 773 -81
rect 781 -101 782 -81
rect 784 -101 785 -81
rect 822 -101 823 -81
rect 825 -101 826 -81
rect 286 -191 287 -171
rect 289 -191 290 -171
rect 155 -239 156 -199
rect 158 -239 159 -199
rect 206 -236 207 -196
rect 209 -236 210 -196
rect 218 -236 219 -196
rect 221 -236 222 -196
rect 252 -236 253 -196
rect 255 -236 256 -196
rect 264 -236 265 -196
rect 267 -236 268 -196
rect 451 -191 452 -171
rect 454 -191 455 -171
rect 320 -239 321 -199
rect 323 -239 324 -199
rect 371 -236 372 -196
rect 374 -236 375 -196
rect 383 -236 384 -196
rect 386 -236 387 -196
rect 417 -236 418 -196
rect 420 -236 421 -196
rect 429 -236 430 -196
rect 432 -236 433 -196
rect 1297 -267 1298 -247
rect 1300 -267 1301 -247
rect 1469 -267 1470 -247
rect 1472 -267 1473 -247
rect 687 -370 688 -350
rect 690 -370 691 -350
rect 699 -370 700 -350
rect 702 -370 703 -350
rect 711 -370 712 -350
rect 714 -370 715 -350
rect 723 -370 724 -350
rect 726 -370 727 -350
rect 760 -370 761 -350
rect 763 -370 764 -350
rect 792 -393 793 -373
rect 795 -393 796 -373
rect 1258 -374 1259 -354
rect 1261 -374 1262 -354
rect 1341 -375 1342 -335
rect 1344 -375 1345 -335
rect 1353 -375 1354 -335
rect 1356 -375 1357 -335
rect 1365 -375 1366 -335
rect 1368 -373 1369 -335
rect 1377 -373 1378 -335
rect 1368 -375 1378 -373
rect 1380 -375 1381 -335
rect 1430 -374 1431 -354
rect 1433 -374 1434 -354
rect 1513 -375 1514 -335
rect 1516 -375 1517 -335
rect 1525 -375 1526 -335
rect 1528 -375 1529 -335
rect 1537 -375 1538 -335
rect 1540 -373 1541 -335
rect 1549 -373 1550 -335
rect 1540 -375 1550 -373
rect 1552 -375 1553 -335
<< pdiffusion >>
rect 706 889 707 929
rect 709 889 710 929
rect 718 889 719 929
rect 721 889 722 929
rect 730 889 731 929
rect 733 889 734 929
rect 742 889 743 929
rect 745 889 746 929
rect 754 889 755 929
rect 757 889 758 929
rect 766 889 767 929
rect 769 889 770 929
rect 778 889 779 929
rect 781 889 782 929
rect 790 889 791 929
rect 793 889 794 929
rect 802 889 803 929
rect 805 889 806 929
rect 814 889 815 929
rect 817 889 818 929
rect 826 889 827 929
rect 829 889 830 929
rect 838 889 839 929
rect 841 889 842 929
rect 850 889 851 929
rect 853 889 854 929
rect 862 889 863 929
rect 865 889 866 929
rect 874 889 875 929
rect 877 889 878 929
rect 912 889 913 929
rect 915 889 916 929
rect 951 889 952 929
rect 954 889 955 929
rect 995 830 996 870
rect 998 830 999 870
rect 1307 654 1308 694
rect 1310 654 1311 694
rect 1351 614 1352 694
rect 1354 614 1355 694
rect 1363 614 1364 694
rect 1366 614 1367 694
rect 1375 614 1376 694
rect 1378 614 1379 694
rect 1387 614 1388 694
rect 1390 614 1391 694
rect 1479 654 1480 694
rect 1482 654 1483 694
rect 1268 547 1269 587
rect 1271 547 1272 587
rect 1523 614 1524 694
rect 1526 614 1527 694
rect 1535 614 1536 694
rect 1538 614 1539 694
rect 1547 614 1548 694
rect 1550 614 1551 694
rect 1559 614 1560 694
rect 1562 614 1563 694
rect 1440 547 1441 587
rect 1443 547 1444 587
rect 696 455 697 495
rect 699 455 700 495
rect 708 455 709 495
rect 711 455 712 495
rect 720 455 721 495
rect 723 455 724 495
rect 732 455 733 495
rect 735 455 736 495
rect 744 455 745 495
rect 747 455 748 495
rect 756 455 757 495
rect 759 455 760 495
rect 768 455 769 495
rect 771 455 772 495
rect 780 455 781 495
rect 783 455 784 495
rect 792 455 793 495
rect 795 455 796 495
rect 804 455 805 495
rect 807 455 808 495
rect 816 455 817 495
rect 819 455 820 495
rect 854 455 855 495
rect 857 455 858 495
rect 893 455 894 495
rect 896 455 897 495
rect 929 385 930 425
rect 932 385 933 425
rect 1302 366 1303 406
rect 1305 366 1306 406
rect 1346 326 1347 406
rect 1349 326 1350 406
rect 1358 326 1359 406
rect 1361 326 1362 406
rect 1370 326 1371 406
rect 1373 326 1374 406
rect 1382 326 1383 406
rect 1385 326 1386 406
rect 1474 366 1475 406
rect 1477 366 1478 406
rect 1263 259 1264 299
rect 1266 259 1267 299
rect 1518 326 1519 406
rect 1521 326 1522 406
rect 1530 326 1531 406
rect 1533 326 1534 406
rect 1542 326 1543 406
rect 1545 326 1546 406
rect 1554 326 1555 406
rect 1557 326 1558 406
rect 1435 259 1436 299
rect 1438 259 1439 299
rect -178 96 -177 176
rect -175 96 -174 176
rect -166 96 -165 176
rect -163 96 -162 176
rect -127 96 -126 176
rect -124 96 -123 176
rect -81 96 -80 176
rect -78 96 -77 176
rect -47 97 -46 137
rect -44 97 -43 137
rect -10 96 -9 176
rect -7 96 -6 176
rect 2 96 3 176
rect 5 96 6 176
rect 41 96 42 176
rect 44 96 45 176
rect 87 96 88 176
rect 90 96 91 176
rect 121 97 122 137
rect 124 97 125 137
rect 156 96 157 176
rect 159 96 160 176
rect 168 96 169 176
rect 171 96 172 176
rect 207 96 208 176
rect 210 96 211 176
rect 253 96 254 176
rect 256 96 257 176
rect 287 97 288 137
rect 290 97 291 137
rect 321 96 322 176
rect 324 96 325 176
rect 333 96 334 176
rect 336 96 337 176
rect 372 96 373 176
rect 375 96 376 176
rect 418 96 419 176
rect 421 96 422 176
rect 452 97 453 137
rect 455 97 456 137
rect 1300 77 1301 117
rect 1303 77 1304 117
rect 697 37 698 77
rect 700 37 701 77
rect 709 37 710 77
rect 712 37 713 77
rect 721 37 722 77
rect 724 37 725 77
rect 733 37 734 77
rect 736 37 737 77
rect 745 37 746 77
rect 748 37 749 77
rect 757 37 758 77
rect 760 37 761 77
rect 769 37 770 77
rect 772 37 773 77
rect 781 37 782 77
rect 784 37 785 77
rect 822 37 823 77
rect 825 37 826 77
rect -179 -155 -178 -75
rect -176 -155 -175 -75
rect -167 -155 -166 -75
rect -164 -155 -163 -75
rect -128 -155 -127 -75
rect -125 -155 -124 -75
rect -82 -155 -81 -75
rect -79 -155 -78 -75
rect -48 -154 -47 -114
rect -45 -154 -44 -114
rect -11 -155 -10 -75
rect -8 -155 -7 -75
rect 1 -155 2 -75
rect 4 -155 5 -75
rect 40 -155 41 -75
rect 43 -155 44 -75
rect 86 -155 87 -75
rect 89 -155 90 -75
rect 120 -154 121 -114
rect 123 -154 124 -114
rect 155 -155 156 -75
rect 158 -155 159 -75
rect 167 -155 168 -75
rect 170 -155 171 -75
rect 206 -155 207 -75
rect 209 -155 210 -75
rect 252 -155 253 -75
rect 255 -155 256 -75
rect 286 -154 287 -114
rect 289 -154 290 -114
rect 320 -155 321 -75
rect 323 -155 324 -75
rect 332 -155 333 -75
rect 335 -155 336 -75
rect 371 -155 372 -75
rect 374 -155 375 -75
rect 417 -155 418 -75
rect 420 -155 421 -75
rect 878 20 879 60
rect 881 20 882 60
rect 1344 37 1345 117
rect 1347 37 1348 117
rect 1356 37 1357 117
rect 1359 37 1360 117
rect 1368 37 1369 117
rect 1371 37 1372 117
rect 1380 37 1381 117
rect 1383 37 1384 117
rect 1472 77 1473 117
rect 1475 77 1476 117
rect 1261 -30 1262 10
rect 1264 -30 1265 10
rect 1516 37 1517 117
rect 1519 37 1520 117
rect 1528 37 1529 117
rect 1531 37 1532 117
rect 1540 37 1541 117
rect 1543 37 1544 117
rect 1552 37 1553 117
rect 1555 37 1556 117
rect 1433 -30 1434 10
rect 1436 -30 1437 10
rect 451 -154 452 -114
rect 454 -154 455 -114
rect 1297 -230 1298 -190
rect 1300 -230 1301 -190
rect 687 -308 688 -268
rect 690 -308 691 -268
rect 699 -308 700 -268
rect 702 -308 703 -268
rect 711 -308 712 -268
rect 714 -308 715 -268
rect 723 -308 724 -268
rect 726 -308 727 -268
rect 760 -308 761 -268
rect 763 -308 764 -268
rect 792 -307 793 -267
rect 795 -307 796 -267
rect 1341 -270 1342 -190
rect 1344 -270 1345 -190
rect 1353 -270 1354 -190
rect 1356 -270 1357 -190
rect 1365 -270 1366 -190
rect 1368 -270 1369 -190
rect 1377 -270 1378 -190
rect 1380 -270 1381 -190
rect 1469 -230 1470 -190
rect 1472 -230 1473 -190
rect 1258 -337 1259 -297
rect 1261 -337 1262 -297
rect 1513 -270 1514 -190
rect 1516 -270 1517 -190
rect 1525 -270 1526 -190
rect 1528 -270 1529 -190
rect 1537 -270 1538 -190
rect 1540 -270 1541 -190
rect 1549 -270 1550 -190
rect 1552 -270 1553 -190
rect 1430 -337 1431 -297
rect 1433 -337 1434 -297
<< ndcontact >>
rect 991 793 995 813
rect 999 793 1003 813
rect 1303 617 1307 637
rect 1311 617 1315 637
rect 1475 617 1479 637
rect 1483 617 1487 637
rect 702 551 706 571
rect 710 551 718 571
rect 722 551 730 571
rect 734 551 742 571
rect 746 551 754 571
rect 758 551 766 571
rect 770 551 778 571
rect 782 551 790 571
rect 794 551 802 571
rect 806 551 814 571
rect 818 551 826 571
rect 830 551 838 571
rect 842 551 850 571
rect 854 551 862 571
rect 866 551 874 571
rect 878 551 882 571
rect 908 551 912 571
rect 916 551 920 571
rect 947 551 951 571
rect 955 551 959 571
rect 1264 510 1268 530
rect 1272 510 1276 530
rect 1347 509 1351 549
rect 1355 509 1363 549
rect 1367 509 1375 549
rect 1379 511 1387 549
rect 1391 509 1395 549
rect 1436 510 1440 530
rect 1444 510 1448 530
rect 1519 509 1523 549
rect 1527 509 1535 549
rect 1539 509 1547 549
rect 1551 511 1559 549
rect 1563 509 1567 549
rect 925 348 929 368
rect 933 348 937 368
rect 1298 329 1302 349
rect 1306 329 1310 349
rect 1470 329 1474 349
rect 1478 329 1482 349
rect 1259 222 1263 242
rect 1267 222 1271 242
rect 1342 221 1346 261
rect 1350 221 1358 261
rect 1362 221 1370 261
rect 1374 223 1382 261
rect 1386 221 1390 261
rect 1431 222 1435 242
rect 1439 222 1443 242
rect 1514 221 1518 261
rect 1522 221 1530 261
rect 1534 221 1542 261
rect 1546 223 1554 261
rect 1558 221 1562 261
rect -51 60 -47 80
rect -43 60 -39 80
rect -182 12 -178 52
rect -174 12 -170 52
rect -131 15 -127 55
rect -123 15 -115 55
rect -111 15 -107 55
rect -85 15 -81 55
rect -77 15 -69 55
rect -65 15 -61 55
rect 117 60 121 80
rect 125 60 129 80
rect -14 12 -10 52
rect -6 12 -2 52
rect 37 15 41 55
rect 45 15 53 55
rect 57 15 61 55
rect 83 15 87 55
rect 91 15 99 55
rect 103 15 107 55
rect 692 164 696 184
rect 700 164 708 184
rect 712 164 720 184
rect 724 164 732 184
rect 736 164 744 184
rect 748 164 756 184
rect 760 164 768 184
rect 772 164 780 184
rect 784 164 792 184
rect 796 164 804 184
rect 808 164 816 184
rect 820 164 824 184
rect 850 164 854 184
rect 858 164 862 184
rect 889 164 893 184
rect 897 164 901 184
rect 283 60 287 80
rect 291 60 295 80
rect 152 12 156 52
rect 160 12 164 52
rect 203 15 207 55
rect 211 15 219 55
rect 223 15 227 55
rect 249 15 253 55
rect 257 15 265 55
rect 269 15 273 55
rect 448 60 452 80
rect 456 60 460 80
rect 317 12 321 52
rect 325 12 329 52
rect 368 15 372 55
rect 376 15 384 55
rect 388 15 392 55
rect 414 15 418 55
rect 422 15 430 55
rect 434 15 438 55
rect -52 -191 -48 -171
rect -44 -191 -40 -171
rect -183 -239 -179 -199
rect -175 -239 -171 -199
rect -132 -236 -128 -196
rect -124 -236 -116 -196
rect -112 -236 -108 -196
rect -86 -236 -82 -196
rect -78 -236 -70 -196
rect -66 -236 -62 -196
rect 116 -191 120 -171
rect 124 -191 128 -171
rect -15 -239 -11 -199
rect -7 -239 -3 -199
rect 36 -236 40 -196
rect 44 -236 52 -196
rect 56 -236 60 -196
rect 82 -236 86 -196
rect 90 -236 98 -196
rect 102 -236 106 -196
rect 1296 40 1300 60
rect 1304 40 1308 60
rect 1468 40 1472 60
rect 1476 40 1480 60
rect 874 -17 878 3
rect 882 -17 886 3
rect 1257 -67 1261 -47
rect 1265 -67 1269 -47
rect 1340 -68 1344 -28
rect 1348 -68 1356 -28
rect 1360 -68 1368 -28
rect 1372 -66 1380 -28
rect 1384 -68 1388 -28
rect 1429 -67 1433 -47
rect 1437 -67 1441 -47
rect 1512 -68 1516 -28
rect 1520 -68 1528 -28
rect 1532 -68 1540 -28
rect 1544 -66 1552 -28
rect 1556 -68 1560 -28
rect 693 -101 697 -81
rect 701 -101 709 -81
rect 713 -101 721 -81
rect 725 -101 733 -81
rect 737 -101 745 -81
rect 749 -101 757 -81
rect 761 -101 769 -81
rect 773 -101 781 -81
rect 785 -101 789 -81
rect 818 -101 822 -81
rect 826 -101 830 -81
rect 282 -191 286 -171
rect 290 -191 294 -171
rect 151 -239 155 -199
rect 159 -239 163 -199
rect 202 -236 206 -196
rect 210 -236 218 -196
rect 222 -236 226 -196
rect 248 -236 252 -196
rect 256 -236 264 -196
rect 268 -236 272 -196
rect 447 -191 451 -171
rect 455 -191 459 -171
rect 316 -239 320 -199
rect 324 -239 328 -199
rect 367 -236 371 -196
rect 375 -236 383 -196
rect 387 -236 391 -196
rect 413 -236 417 -196
rect 421 -236 429 -196
rect 433 -236 437 -196
rect 1293 -267 1297 -247
rect 1301 -267 1305 -247
rect 1465 -267 1469 -247
rect 1473 -267 1477 -247
rect 683 -370 687 -350
rect 691 -370 699 -350
rect 703 -370 711 -350
rect 715 -370 723 -350
rect 727 -370 731 -350
rect 756 -370 760 -350
rect 764 -370 768 -350
rect 788 -393 792 -373
rect 796 -393 800 -373
rect 1254 -374 1258 -354
rect 1262 -374 1266 -354
rect 1337 -375 1341 -335
rect 1345 -375 1353 -335
rect 1357 -375 1365 -335
rect 1369 -373 1377 -335
rect 1381 -375 1385 -335
rect 1426 -374 1430 -354
rect 1434 -374 1438 -354
rect 1509 -375 1513 -335
rect 1517 -375 1525 -335
rect 1529 -375 1537 -335
rect 1541 -373 1549 -335
rect 1553 -375 1557 -335
<< pdcontact >>
rect 702 889 706 929
rect 710 889 718 929
rect 722 889 730 929
rect 734 889 742 929
rect 746 889 754 929
rect 758 889 766 929
rect 770 889 778 929
rect 782 889 790 929
rect 794 889 802 929
rect 806 889 814 929
rect 818 889 826 929
rect 830 889 838 929
rect 842 889 850 929
rect 854 889 862 929
rect 866 889 874 929
rect 878 889 882 929
rect 908 889 912 929
rect 916 889 920 929
rect 947 889 951 929
rect 955 889 959 929
rect 991 830 995 870
rect 999 830 1003 870
rect 1303 654 1307 694
rect 1311 654 1315 694
rect 1347 614 1351 694
rect 1355 614 1363 694
rect 1367 614 1375 694
rect 1379 614 1387 694
rect 1391 614 1395 694
rect 1475 654 1479 694
rect 1483 654 1487 694
rect 1264 547 1268 587
rect 1272 547 1276 587
rect 1519 614 1523 694
rect 1527 614 1535 694
rect 1539 614 1547 694
rect 1551 614 1559 694
rect 1563 614 1567 694
rect 1436 547 1440 587
rect 1444 547 1448 587
rect 692 455 696 495
rect 700 455 708 495
rect 712 455 720 495
rect 724 455 732 495
rect 736 455 744 495
rect 748 455 756 495
rect 760 455 768 495
rect 772 455 780 495
rect 784 455 792 495
rect 796 455 804 495
rect 808 455 816 495
rect 820 455 824 495
rect 850 455 854 495
rect 858 455 862 495
rect 889 455 893 495
rect 897 455 901 495
rect 925 385 929 425
rect 933 385 937 425
rect 1298 366 1302 406
rect 1306 366 1310 406
rect 1342 326 1346 406
rect 1350 326 1358 406
rect 1362 326 1370 406
rect 1374 326 1382 406
rect 1386 326 1390 406
rect 1470 366 1474 406
rect 1478 366 1482 406
rect 1259 259 1263 299
rect 1267 259 1271 299
rect 1514 326 1518 406
rect 1522 326 1530 406
rect 1534 326 1542 406
rect 1546 326 1554 406
rect 1558 326 1562 406
rect 1431 259 1435 299
rect 1439 259 1443 299
rect -182 96 -178 176
rect -174 96 -166 176
rect -162 96 -158 176
rect -131 96 -127 176
rect -123 96 -119 176
rect -85 96 -81 176
rect -77 96 -73 176
rect -51 97 -47 137
rect -43 97 -39 137
rect -14 96 -10 176
rect -6 96 2 176
rect 6 96 10 176
rect 37 96 41 176
rect 45 96 49 176
rect 83 96 87 176
rect 91 96 95 176
rect 117 97 121 137
rect 125 97 129 137
rect 152 96 156 176
rect 160 96 168 176
rect 172 96 176 176
rect 203 96 207 176
rect 211 96 215 176
rect 249 96 253 176
rect 257 96 261 176
rect 283 97 287 137
rect 291 97 295 137
rect 317 96 321 176
rect 325 96 333 176
rect 337 96 341 176
rect 368 96 372 176
rect 376 96 380 176
rect 414 96 418 176
rect 422 96 426 176
rect 448 97 452 137
rect 456 97 460 137
rect 1296 77 1300 117
rect 1304 77 1308 117
rect 693 37 697 77
rect 701 37 709 77
rect 713 37 721 77
rect 725 37 733 77
rect 737 37 745 77
rect 749 37 757 77
rect 761 37 769 77
rect 773 37 781 77
rect 785 37 789 77
rect 818 37 822 77
rect 826 37 830 77
rect -183 -155 -179 -75
rect -175 -155 -167 -75
rect -163 -155 -159 -75
rect -132 -155 -128 -75
rect -124 -155 -120 -75
rect -86 -155 -82 -75
rect -78 -155 -74 -75
rect -52 -154 -48 -114
rect -44 -154 -40 -114
rect -15 -155 -11 -75
rect -7 -155 1 -75
rect 5 -155 9 -75
rect 36 -155 40 -75
rect 44 -155 48 -75
rect 82 -155 86 -75
rect 90 -155 94 -75
rect 116 -154 120 -114
rect 124 -154 128 -114
rect 151 -155 155 -75
rect 159 -155 167 -75
rect 171 -155 175 -75
rect 202 -155 206 -75
rect 210 -155 214 -75
rect 248 -155 252 -75
rect 256 -155 260 -75
rect 282 -154 286 -114
rect 290 -154 294 -114
rect 316 -155 320 -75
rect 324 -155 332 -75
rect 336 -155 340 -75
rect 367 -155 371 -75
rect 375 -155 379 -75
rect 413 -155 417 -75
rect 421 -155 425 -75
rect 874 20 878 60
rect 882 20 886 60
rect 1340 37 1344 117
rect 1348 37 1356 117
rect 1360 37 1368 117
rect 1372 37 1380 117
rect 1384 37 1388 117
rect 1468 77 1472 117
rect 1476 77 1480 117
rect 1257 -30 1261 10
rect 1265 -30 1269 10
rect 1512 37 1516 117
rect 1520 37 1528 117
rect 1532 37 1540 117
rect 1544 37 1552 117
rect 1556 37 1560 117
rect 1429 -30 1433 10
rect 1437 -30 1441 10
rect 447 -154 451 -114
rect 455 -154 459 -114
rect 1293 -230 1297 -190
rect 1301 -230 1305 -190
rect 683 -308 687 -268
rect 691 -308 699 -268
rect 703 -308 711 -268
rect 715 -308 723 -268
rect 727 -308 731 -268
rect 756 -308 760 -268
rect 764 -308 768 -268
rect 788 -307 792 -267
rect 796 -307 800 -267
rect 1337 -270 1341 -190
rect 1345 -270 1353 -190
rect 1357 -270 1365 -190
rect 1369 -270 1377 -190
rect 1381 -270 1385 -190
rect 1465 -230 1469 -190
rect 1473 -230 1477 -190
rect 1254 -337 1258 -297
rect 1262 -337 1266 -297
rect 1509 -270 1513 -190
rect 1517 -270 1525 -190
rect 1529 -270 1537 -190
rect 1541 -270 1549 -190
rect 1553 -270 1557 -190
rect 1426 -337 1430 -297
rect 1434 -337 1438 -297
<< polysilicon >>
rect 707 929 709 932
rect 719 929 721 933
rect 731 929 733 932
rect 743 929 745 932
rect 755 929 757 932
rect 767 929 769 932
rect 779 929 781 932
rect 791 929 793 932
rect 803 929 805 932
rect 815 929 817 932
rect 827 929 829 932
rect 839 929 841 932
rect 851 929 853 932
rect 863 929 865 932
rect 875 929 877 932
rect 913 929 915 932
rect 952 929 954 932
rect 707 571 709 889
rect 719 571 721 889
rect 731 571 733 889
rect 743 571 745 889
rect 755 571 757 889
rect 767 571 769 889
rect 779 571 781 889
rect 791 571 793 889
rect 803 571 805 889
rect 815 571 817 889
rect 827 571 829 889
rect 839 571 841 889
rect 851 571 853 889
rect 863 571 865 889
rect 875 571 877 889
rect 913 571 915 889
rect 952 571 954 889
rect 996 870 998 876
rect 996 813 998 830
rect 996 789 998 793
rect 1308 694 1310 700
rect 1352 694 1354 698
rect 1364 694 1366 698
rect 1376 694 1378 698
rect 1388 694 1390 698
rect 1480 694 1482 700
rect 1524 694 1526 698
rect 1536 694 1538 698
rect 1548 694 1550 698
rect 1560 694 1562 698
rect 1308 637 1310 654
rect 1308 613 1310 617
rect 1480 637 1482 654
rect 1269 587 1271 593
rect 707 547 709 551
rect 719 548 721 551
rect 731 548 733 551
rect 743 547 745 551
rect 755 546 757 551
rect 767 546 769 551
rect 779 546 781 551
rect 791 547 793 551
rect 803 547 805 551
rect 815 546 817 551
rect 827 546 829 551
rect 839 546 841 551
rect 851 547 853 551
rect 863 547 865 551
rect 875 547 877 551
rect 913 547 915 551
rect 952 547 954 551
rect 1352 549 1354 614
rect 1364 549 1366 614
rect 1376 549 1378 614
rect 1388 549 1390 614
rect 1480 613 1482 617
rect 1441 587 1443 593
rect 1269 530 1271 547
rect 1269 506 1271 510
rect 1524 549 1526 614
rect 1536 549 1538 614
rect 1548 549 1550 614
rect 1560 549 1562 614
rect 1441 530 1443 547
rect 1352 505 1354 509
rect 1364 505 1366 509
rect 1376 504 1378 509
rect 1388 504 1390 509
rect 1441 506 1443 510
rect 1524 505 1526 509
rect 1536 505 1538 509
rect 1548 504 1550 509
rect 1560 504 1562 509
rect 697 495 699 498
rect 709 495 711 498
rect 721 495 723 498
rect 733 495 735 498
rect 745 495 747 498
rect 757 495 759 498
rect 769 495 771 498
rect 781 495 783 498
rect 793 495 795 498
rect 805 495 807 498
rect 817 495 819 498
rect 855 495 857 498
rect 894 495 896 498
rect 697 184 699 455
rect 709 184 711 455
rect 721 184 723 455
rect 733 184 735 455
rect 745 184 747 455
rect 757 184 759 455
rect 769 184 771 455
rect 781 184 783 455
rect 793 184 795 455
rect 805 184 807 455
rect 817 184 819 455
rect 855 184 857 455
rect 894 184 896 455
rect 930 425 932 431
rect 1303 406 1305 412
rect 1347 406 1349 410
rect 1359 406 1361 410
rect 1371 406 1373 410
rect 1383 406 1385 410
rect 1475 406 1477 412
rect 1519 406 1521 410
rect 1531 406 1533 410
rect 1543 406 1545 410
rect 1555 406 1557 410
rect 930 368 932 385
rect 1303 349 1305 366
rect 930 344 932 348
rect 1303 325 1305 329
rect 1475 349 1477 366
rect 1264 299 1266 305
rect 1347 261 1349 326
rect 1359 261 1361 326
rect 1371 261 1373 326
rect 1383 261 1385 326
rect 1475 325 1477 329
rect 1436 299 1438 305
rect 1264 242 1266 259
rect 1264 218 1266 222
rect 1519 261 1521 326
rect 1531 261 1533 326
rect 1543 261 1545 326
rect 1555 261 1557 326
rect 1436 242 1438 259
rect 1347 217 1349 221
rect 1359 217 1361 221
rect 1371 216 1373 221
rect 1383 216 1385 221
rect 1436 218 1438 222
rect 1519 217 1521 221
rect 1531 217 1533 221
rect 1543 216 1545 221
rect 1555 216 1557 221
rect -177 176 -175 180
rect -165 176 -163 180
rect -126 176 -124 180
rect -80 176 -78 180
rect -9 176 -7 180
rect 3 176 5 180
rect 42 176 44 180
rect 88 176 90 180
rect 157 176 159 180
rect 169 176 171 180
rect 208 176 210 180
rect 254 176 256 180
rect 322 176 324 180
rect 334 176 336 180
rect 373 176 375 180
rect 419 176 421 180
rect -46 137 -44 143
rect -177 52 -175 96
rect -165 72 -163 96
rect -126 79 -124 96
rect -80 79 -78 96
rect -46 80 -44 97
rect 122 137 124 143
rect -126 55 -124 66
rect -114 55 -112 67
rect -80 55 -78 66
rect -68 55 -66 67
rect -46 56 -44 60
rect -9 52 -7 96
rect 3 72 5 96
rect 42 79 44 96
rect 88 79 90 96
rect 122 80 124 97
rect 288 137 290 143
rect 42 55 44 66
rect 54 55 56 67
rect 88 55 90 66
rect 100 55 102 67
rect 122 56 124 60
rect -177 6 -175 12
rect -126 11 -124 15
rect -114 12 -112 15
rect -80 11 -78 15
rect -68 12 -66 15
rect 157 52 159 96
rect 169 72 171 96
rect 208 79 210 96
rect 254 79 256 96
rect 288 80 290 97
rect 697 159 699 164
rect 709 159 711 164
rect 721 159 723 164
rect 733 160 735 164
rect 745 160 747 164
rect 757 159 759 164
rect 769 159 771 164
rect 781 159 783 164
rect 793 160 795 164
rect 805 160 807 164
rect 817 160 819 164
rect 855 160 857 164
rect 894 160 896 164
rect 453 137 455 143
rect 1301 117 1303 123
rect 1345 117 1347 121
rect 1357 117 1359 121
rect 1369 117 1371 121
rect 1381 117 1383 121
rect 1473 117 1475 123
rect 1517 117 1519 121
rect 1529 117 1531 121
rect 1541 117 1543 121
rect 1553 117 1555 121
rect 208 55 210 66
rect 220 55 222 67
rect 254 55 256 66
rect 266 55 268 67
rect 288 56 290 60
rect -9 6 -7 12
rect 42 11 44 15
rect 54 12 56 15
rect 88 11 90 15
rect 100 12 102 15
rect 322 52 324 96
rect 334 72 336 96
rect 373 79 375 96
rect 419 79 421 96
rect 453 80 455 97
rect 373 55 375 66
rect 385 55 387 67
rect 419 55 421 66
rect 431 55 433 67
rect 698 77 700 80
rect 710 77 712 80
rect 722 77 724 80
rect 734 77 736 80
rect 746 77 748 80
rect 758 77 760 80
rect 770 77 772 80
rect 782 77 784 80
rect 823 77 825 81
rect 453 56 455 60
rect 157 6 159 12
rect 208 11 210 15
rect 220 12 222 15
rect 254 11 256 15
rect 266 12 268 15
rect 879 60 881 66
rect 1301 60 1303 77
rect 322 6 324 12
rect 373 11 375 15
rect 385 12 387 15
rect 419 11 421 15
rect 431 12 433 15
rect -178 -75 -176 -71
rect -166 -75 -164 -71
rect -127 -75 -125 -71
rect -81 -75 -79 -71
rect -10 -75 -8 -71
rect 2 -75 4 -71
rect 41 -75 43 -71
rect 87 -75 89 -71
rect 156 -75 158 -71
rect 168 -75 170 -71
rect 207 -75 209 -71
rect 253 -75 255 -71
rect 321 -75 323 -71
rect 333 -75 335 -71
rect 372 -75 374 -71
rect 418 -75 420 -71
rect -47 -114 -45 -108
rect -178 -199 -176 -155
rect -166 -179 -164 -155
rect -127 -172 -125 -155
rect -81 -172 -79 -155
rect -47 -171 -45 -154
rect 121 -114 123 -108
rect -127 -196 -125 -185
rect -115 -196 -113 -184
rect -81 -196 -79 -185
rect -69 -196 -67 -184
rect -47 -195 -45 -191
rect -10 -199 -8 -155
rect 2 -179 4 -155
rect 41 -172 43 -155
rect 87 -172 89 -155
rect 121 -171 123 -154
rect 287 -114 289 -108
rect 41 -196 43 -185
rect 53 -196 55 -184
rect 87 -196 89 -185
rect 99 -196 101 -184
rect 121 -195 123 -191
rect -178 -245 -176 -239
rect -127 -240 -125 -236
rect -115 -239 -113 -236
rect -81 -240 -79 -236
rect -69 -239 -67 -236
rect 156 -199 158 -155
rect 168 -179 170 -155
rect 207 -172 209 -155
rect 253 -172 255 -155
rect 287 -171 289 -154
rect 698 -81 700 37
rect 710 -81 712 37
rect 722 -81 724 37
rect 734 -81 736 37
rect 746 -81 748 37
rect 758 -81 760 37
rect 770 -81 772 37
rect 782 -81 784 37
rect 823 -81 825 37
rect 1301 36 1303 40
rect 1473 60 1475 77
rect 879 3 881 20
rect 1262 10 1264 16
rect 879 -21 881 -17
rect 1345 -28 1347 37
rect 1357 -28 1359 37
rect 1369 -28 1371 37
rect 1381 -28 1383 37
rect 1473 36 1475 40
rect 1434 10 1436 16
rect 1262 -47 1264 -30
rect 1262 -71 1264 -67
rect 1517 -28 1519 37
rect 1529 -28 1531 37
rect 1541 -28 1543 37
rect 1553 -28 1555 37
rect 1434 -47 1436 -30
rect 1345 -72 1347 -68
rect 1357 -72 1359 -68
rect 1369 -73 1371 -68
rect 1381 -73 1383 -68
rect 1434 -71 1436 -67
rect 1517 -72 1519 -68
rect 1529 -72 1531 -68
rect 1541 -73 1543 -68
rect 1553 -73 1555 -68
rect 698 -105 700 -101
rect 710 -105 712 -101
rect 722 -105 724 -101
rect 734 -105 736 -101
rect 746 -105 748 -101
rect 758 -105 760 -101
rect 770 -105 772 -101
rect 782 -105 784 -101
rect 823 -105 825 -101
rect 452 -114 454 -108
rect 207 -196 209 -185
rect 219 -196 221 -184
rect 253 -196 255 -185
rect 265 -196 267 -184
rect 287 -195 289 -191
rect -10 -245 -8 -239
rect 41 -240 43 -236
rect 53 -239 55 -236
rect 87 -240 89 -236
rect 99 -239 101 -236
rect 321 -199 323 -155
rect 333 -179 335 -155
rect 372 -172 374 -155
rect 418 -172 420 -155
rect 452 -171 454 -154
rect 372 -196 374 -185
rect 384 -196 386 -184
rect 418 -196 420 -185
rect 430 -196 432 -184
rect 1298 -190 1300 -184
rect 1342 -190 1344 -186
rect 1354 -190 1356 -186
rect 1366 -190 1368 -186
rect 1378 -190 1380 -186
rect 1470 -190 1472 -184
rect 1514 -190 1516 -186
rect 1526 -190 1528 -186
rect 1538 -190 1540 -186
rect 1550 -190 1552 -186
rect 452 -195 454 -191
rect 156 -245 158 -239
rect 207 -240 209 -236
rect 219 -239 221 -236
rect 253 -240 255 -236
rect 265 -239 267 -236
rect 321 -245 323 -239
rect 372 -240 374 -236
rect 384 -239 386 -236
rect 418 -240 420 -236
rect 430 -239 432 -236
rect 1298 -247 1300 -230
rect 688 -268 690 -265
rect 700 -268 702 -265
rect 712 -268 714 -265
rect 724 -268 726 -265
rect 761 -268 763 -265
rect 793 -267 795 -261
rect 1298 -271 1300 -267
rect 1470 -247 1472 -230
rect 1259 -297 1261 -291
rect 688 -350 690 -308
rect 700 -350 702 -308
rect 712 -350 714 -308
rect 724 -350 726 -308
rect 761 -350 763 -308
rect 688 -375 690 -370
rect 700 -375 702 -370
rect 712 -374 714 -370
rect 724 -374 726 -370
rect 761 -374 763 -370
rect 793 -373 795 -307
rect 1342 -335 1344 -270
rect 1354 -335 1356 -270
rect 1366 -335 1368 -270
rect 1378 -335 1380 -270
rect 1470 -271 1472 -267
rect 1431 -297 1433 -291
rect 1259 -354 1261 -337
rect 1259 -378 1261 -374
rect 1514 -335 1516 -270
rect 1526 -335 1528 -270
rect 1538 -335 1540 -270
rect 1550 -335 1552 -270
rect 1431 -354 1433 -337
rect 1342 -379 1344 -375
rect 1354 -379 1356 -375
rect 1366 -380 1368 -375
rect 1378 -380 1380 -375
rect 1431 -378 1433 -374
rect 1514 -379 1516 -375
rect 1526 -379 1528 -375
rect 1538 -380 1540 -375
rect 1550 -380 1552 -375
rect 793 -397 795 -393
<< polycontact >>
rect 702 796 707 802
rect 714 785 719 790
rect 733 777 738 782
rect 738 768 743 773
rect 750 758 755 764
rect 762 749 767 754
rect 774 741 779 746
rect 786 732 791 737
rect 798 723 803 728
rect 810 714 815 719
rect 822 705 827 710
rect 834 696 839 701
rect 846 687 851 692
rect 858 678 863 683
rect 870 669 875 674
rect 908 660 913 665
rect 947 651 952 656
rect 991 817 996 821
rect 1303 641 1308 645
rect 1475 641 1480 645
rect 1346 591 1352 595
rect 1359 583 1364 587
rect 1371 573 1376 577
rect 1384 563 1388 567
rect 1518 591 1524 595
rect 1264 534 1269 538
rect 1531 583 1536 587
rect 1543 573 1548 577
rect 1556 563 1560 567
rect 1436 534 1441 538
rect 693 360 697 364
rect 705 351 709 355
rect 723 343 727 347
rect 729 335 733 339
rect 741 325 745 329
rect 753 317 757 321
rect 765 309 769 313
rect 777 300 781 305
rect 789 290 793 295
rect 801 278 805 283
rect 813 268 817 273
rect 851 258 855 263
rect 890 249 894 254
rect 925 372 930 376
rect 1298 353 1303 357
rect 1470 353 1475 357
rect 1341 303 1347 307
rect 1354 295 1359 299
rect 1366 285 1371 289
rect 1379 275 1383 279
rect 1513 303 1519 307
rect 1259 246 1264 250
rect 1526 295 1531 299
rect 1538 285 1543 289
rect 1551 275 1555 279
rect 1431 246 1436 250
rect -183 67 -177 72
rect -51 83 -46 87
rect -163 75 -157 79
rect -128 75 -122 79
rect -82 75 -76 79
rect -127 66 -123 70
rect -115 67 -111 72
rect -81 66 -77 70
rect -69 67 -65 72
rect -15 67 -9 72
rect 117 83 122 87
rect 5 75 11 79
rect 40 75 46 79
rect 86 75 92 79
rect 41 66 45 70
rect 53 67 57 72
rect 87 66 91 70
rect 99 67 103 72
rect 151 67 157 72
rect 283 83 288 87
rect 171 75 177 79
rect 206 75 212 79
rect 252 75 258 79
rect 207 66 211 70
rect 219 67 223 72
rect 253 66 257 70
rect 265 67 269 72
rect 316 67 322 72
rect 448 83 453 87
rect 336 75 342 79
rect 371 75 377 79
rect 417 75 423 79
rect 372 66 376 70
rect 384 67 388 72
rect 418 66 422 70
rect 430 67 434 72
rect 1296 64 1301 68
rect 694 -1 698 3
rect -184 -184 -178 -179
rect -52 -168 -47 -164
rect -164 -176 -158 -172
rect -129 -176 -123 -172
rect -83 -176 -77 -172
rect -128 -185 -124 -181
rect -116 -184 -112 -179
rect -82 -185 -78 -181
rect -70 -184 -66 -179
rect -16 -184 -10 -179
rect 116 -168 121 -164
rect 4 -176 10 -172
rect 39 -176 45 -172
rect 85 -176 91 -172
rect 40 -185 44 -181
rect 52 -184 56 -179
rect 86 -185 90 -181
rect 98 -184 102 -179
rect 150 -184 156 -179
rect 282 -168 287 -164
rect 706 -10 710 -6
rect 724 -18 729 -14
rect 729 -26 734 -22
rect 742 -35 746 -31
rect 754 -43 758 -39
rect 766 -52 770 -48
rect 778 -59 782 -55
rect 1468 64 1473 68
rect 874 7 879 11
rect 1339 14 1345 18
rect 1352 6 1357 10
rect 1364 -4 1369 0
rect 1377 -14 1381 -10
rect 1511 14 1517 18
rect 1257 -43 1262 -39
rect 1524 6 1529 10
rect 1536 -4 1541 0
rect 1549 -14 1553 -10
rect 1429 -43 1434 -39
rect 170 -176 176 -172
rect 205 -176 211 -172
rect 251 -176 257 -172
rect 206 -185 210 -181
rect 218 -184 222 -179
rect 252 -185 256 -181
rect 264 -184 268 -179
rect 315 -184 321 -179
rect 447 -168 452 -164
rect 335 -176 341 -172
rect 370 -176 376 -172
rect 416 -176 422 -172
rect 371 -185 375 -181
rect 383 -184 387 -179
rect 417 -185 421 -181
rect 429 -184 433 -179
rect 1293 -243 1298 -239
rect 687 -265 691 -261
rect 699 -265 703 -261
rect 711 -265 715 -261
rect 723 -265 727 -261
rect 760 -265 764 -261
rect 1465 -243 1470 -239
rect 1336 -293 1342 -289
rect 788 -347 793 -343
rect 1349 -301 1354 -297
rect 1361 -311 1366 -307
rect 1374 -321 1378 -317
rect 1508 -293 1514 -289
rect 1254 -350 1259 -346
rect 1521 -301 1526 -297
rect 1533 -311 1538 -307
rect 1546 -321 1550 -317
rect 1426 -350 1431 -346
<< metal1 >>
rect 525 942 1028 946
rect 525 517 529 942
rect 702 929 706 942
rect 760 929 765 942
rect 844 929 849 942
rect 991 941 1028 942
rect 724 822 728 889
rect 736 833 741 889
rect 784 848 789 889
rect 796 871 801 889
rect 808 848 813 889
rect 819 868 824 889
rect 856 877 861 889
rect 867 887 872 889
rect 878 887 882 889
rect 909 877 912 889
rect 856 872 912 877
rect 916 868 920 889
rect 819 863 867 868
rect 872 863 920 868
rect 784 842 878 848
rect 736 829 795 833
rect 948 833 951 889
rect 802 829 951 833
rect 955 821 959 889
rect 991 870 994 941
rect 999 821 1003 830
rect 729 817 991 821
rect 999 817 1016 821
rect 724 808 728 813
rect 600 797 681 802
rect 595 796 681 797
rect 691 796 702 802
rect 662 785 714 790
rect 702 781 707 785
rect 702 777 733 781
rect 738 777 739 781
rect 702 776 739 777
rect 651 768 711 773
rect 717 768 738 773
rect 583 763 735 764
rect 588 758 735 763
rect 741 758 750 764
rect 574 749 698 754
rect 704 749 762 754
rect 641 741 747 746
rect 752 741 774 746
rect 717 732 786 737
rect 741 723 798 728
rect 752 714 810 719
rect 631 705 808 710
rect 813 705 822 710
rect 563 696 820 701
rect 826 696 834 701
rect 665 687 667 692
rect 673 687 846 692
rect 826 678 858 683
rect 704 669 870 674
rect 813 660 908 665
rect 680 651 681 656
rect 691 651 947 656
rect 736 639 794 645
rect 724 571 728 576
rect 736 571 741 639
rect 801 639 951 645
rect 784 626 878 631
rect 784 571 788 626
rect 795 571 800 583
rect 808 571 812 626
rect 819 596 867 603
rect 873 596 920 603
rect 819 571 823 596
rect 856 582 912 587
rect 856 571 860 582
rect 878 571 882 572
rect 908 571 912 582
rect 916 571 920 596
rect 947 571 951 639
rect 955 571 959 817
rect 999 813 1003 817
rect 702 541 706 551
rect 760 541 764 551
rect 844 541 848 551
rect 991 541 995 793
rect 701 536 995 541
rect 525 513 928 517
rect 525 190 529 513
rect 692 495 696 513
rect 750 495 754 513
rect 820 495 824 513
rect 714 376 718 455
rect 726 403 730 455
rect 774 426 778 455
rect 786 403 790 455
rect 798 426 802 455
rect 810 437 814 455
rect 851 437 854 455
rect 810 434 854 437
rect 858 427 862 455
rect 890 403 893 455
rect 726 399 893 403
rect 897 376 901 455
rect 925 425 928 513
rect 933 376 937 385
rect 719 372 925 376
rect 933 372 945 376
rect 719 371 901 372
rect 589 360 686 364
rect 692 360 693 364
rect 652 351 705 355
rect 692 347 696 351
rect 692 343 723 347
rect 727 343 729 347
rect 642 335 701 339
rect 706 335 729 339
rect 576 325 725 329
rect 731 325 741 329
rect 564 317 737 321
rect 742 317 753 321
rect 632 309 749 313
rect 755 309 765 313
rect 706 300 777 305
rect 731 290 789 295
rect 737 278 738 283
rect 743 278 801 283
rect 676 268 813 273
rect 755 258 851 263
rect 692 249 890 254
rect 726 233 893 237
rect -208 182 529 190
rect 714 184 718 227
rect 726 184 730 233
rect 774 184 777 204
rect 787 184 791 233
rect 799 184 802 205
rect 810 190 853 195
rect 810 184 813 190
rect 850 184 853 190
rect 858 184 861 205
rect 889 184 893 233
rect -208 -61 -197 182
rect -182 176 -178 182
rect -131 176 -127 182
rect -85 176 -81 182
rect -51 181 529 182
rect -51 137 -47 181
rect -14 176 -10 181
rect 37 176 41 181
rect 83 176 87 181
rect -162 86 -158 96
rect -174 82 -158 86
rect -123 87 -119 96
rect -136 83 -98 87
rect -77 87 -73 96
rect -43 88 -39 97
rect 117 137 121 181
rect 152 176 156 181
rect 203 176 207 181
rect 249 176 253 181
rect -90 83 -51 87
rect -43 84 -33 88
rect -27 84 -25 88
rect 6 86 10 96
rect -188 67 -183 72
rect -174 70 -170 82
rect -157 75 -151 79
rect -101 79 -98 83
rect -43 80 -39 84
rect -146 75 -128 79
rect -122 75 -104 79
rect -101 75 -82 79
rect -76 75 -65 79
rect -115 72 -111 75
rect -174 66 -127 70
rect -108 70 -104 75
rect -69 72 -65 75
rect -108 66 -81 70
rect -174 52 -170 66
rect -6 82 10 86
rect 45 87 49 96
rect 32 83 70 87
rect 91 87 95 96
rect 125 88 129 97
rect 283 137 287 181
rect 317 176 321 181
rect 368 176 372 181
rect 414 176 418 181
rect 78 83 117 87
rect 125 84 137 88
rect -20 67 -15 72
rect -6 70 -2 82
rect 11 75 17 79
rect 67 79 70 83
rect 125 80 129 84
rect 142 84 143 88
rect 172 86 176 96
rect 22 75 40 79
rect 46 75 64 79
rect 67 75 86 79
rect 92 75 103 79
rect 53 72 57 75
rect -6 66 41 70
rect 60 70 64 75
rect 99 72 103 75
rect 60 66 87 70
rect -182 6 -178 12
rect -111 6 -107 15
rect -65 6 -61 15
rect -51 6 -46 60
rect -6 52 -2 66
rect 160 82 176 86
rect 211 87 215 96
rect 198 83 236 87
rect 257 87 261 96
rect 291 88 295 97
rect 448 137 452 181
rect 244 83 283 87
rect 291 84 301 88
rect 146 67 151 72
rect 160 70 164 82
rect 177 75 183 79
rect 233 79 236 83
rect 291 80 295 84
rect 337 86 341 96
rect 188 75 206 79
rect 212 75 230 79
rect 233 75 252 79
rect 258 75 269 79
rect 219 72 223 75
rect 160 66 207 70
rect 226 70 230 75
rect 265 72 269 75
rect 226 66 253 70
rect -14 6 -10 12
rect 57 6 61 15
rect 103 6 107 15
rect 117 6 122 60
rect 160 52 164 66
rect 325 82 341 86
rect 376 87 380 96
rect 363 83 401 87
rect 422 87 426 96
rect 456 88 460 97
rect 525 107 529 181
rect 897 184 901 371
rect 933 368 937 372
rect 692 143 696 164
rect 750 143 754 164
rect 820 143 824 164
rect 925 143 929 348
rect 991 143 995 536
rect 1024 704 1028 941
rect 1089 724 1409 732
rect 1024 700 1573 704
rect 1024 699 1268 700
rect 1024 417 1028 699
rect 1229 641 1256 645
rect 1264 587 1268 699
rect 1303 694 1307 700
rect 1367 694 1375 700
rect 1311 645 1315 654
rect 1282 641 1303 645
rect 1311 641 1326 645
rect 1283 579 1288 641
rect 1311 637 1315 641
rect 1154 534 1252 538
rect 1272 538 1276 547
rect 1257 534 1264 538
rect 1272 534 1291 538
rect 1272 530 1276 534
rect 1264 502 1268 510
rect 1303 502 1307 617
rect 1322 595 1326 641
rect 1419 641 1428 645
rect 1347 606 1351 614
rect 1391 606 1395 614
rect 1347 601 1412 606
rect 1322 591 1346 595
rect 1330 583 1359 587
rect 1329 573 1371 577
rect 1322 563 1384 567
rect 1322 539 1327 563
rect 1347 553 1395 558
rect 1347 549 1351 553
rect 1391 549 1395 553
rect 1379 509 1387 511
rect 1357 502 1361 509
rect 1264 498 1361 502
rect 1381 502 1385 509
rect 1399 502 1403 601
rect 1407 538 1412 601
rect 1436 587 1440 700
rect 1475 694 1479 700
rect 1539 694 1547 700
rect 1483 645 1487 654
rect 1454 641 1475 645
rect 1483 641 1498 645
rect 1455 579 1460 641
rect 1483 637 1487 641
rect 1407 534 1424 538
rect 1444 538 1448 547
rect 1429 534 1436 538
rect 1444 534 1463 538
rect 1444 530 1448 534
rect 1381 498 1403 502
rect 1436 502 1440 510
rect 1475 502 1479 617
rect 1494 595 1498 641
rect 1519 606 1523 614
rect 1563 606 1567 614
rect 1519 601 1581 606
rect 1494 591 1518 595
rect 1502 583 1531 587
rect 1501 573 1543 577
rect 1494 563 1556 567
rect 1494 539 1499 563
rect 1519 553 1567 558
rect 1519 549 1523 553
rect 1563 549 1567 553
rect 1551 509 1559 511
rect 1529 502 1533 509
rect 1436 498 1533 502
rect 1553 502 1557 509
rect 1571 502 1575 601
rect 1553 498 1575 502
rect 1356 491 1361 498
rect 1436 492 1440 498
rect 1436 491 1602 492
rect 1356 485 1602 491
rect 1078 436 1404 444
rect 1023 416 1259 417
rect 1023 412 1568 416
rect 1023 411 1263 412
rect 692 138 995 143
rect 525 103 877 107
rect 409 83 448 87
rect 456 84 470 88
rect 311 67 316 72
rect 325 70 329 82
rect 342 75 348 79
rect 398 79 401 83
rect 456 80 460 84
rect 353 75 371 79
rect 377 75 395 79
rect 398 75 417 79
rect 423 75 434 79
rect 384 72 388 75
rect 325 66 372 70
rect 391 70 395 75
rect 430 72 434 75
rect 391 66 418 70
rect 152 6 156 12
rect 223 6 227 15
rect 269 6 273 15
rect 283 6 288 60
rect 325 52 329 66
rect 317 6 321 12
rect 388 6 392 15
rect 434 6 438 15
rect 448 6 453 60
rect -186 1 502 6
rect -208 -69 451 -61
rect -183 -75 -179 -69
rect -132 -75 -128 -69
rect -86 -75 -82 -69
rect -52 -70 451 -69
rect -52 -114 -48 -70
rect -15 -75 -11 -70
rect 36 -75 40 -70
rect 82 -75 86 -70
rect -163 -165 -159 -155
rect -175 -169 -159 -165
rect -124 -164 -120 -155
rect -137 -168 -99 -164
rect -78 -164 -74 -155
rect -44 -163 -40 -154
rect 116 -114 120 -70
rect 151 -75 155 -70
rect 202 -75 206 -70
rect 248 -75 252 -70
rect -91 -168 -52 -164
rect -44 -167 -34 -163
rect -28 -167 -26 -163
rect 5 -165 9 -155
rect -189 -184 -184 -179
rect -175 -181 -171 -169
rect -158 -176 -152 -172
rect -102 -172 -99 -168
rect -44 -171 -40 -167
rect -147 -176 -129 -172
rect -123 -176 -105 -172
rect -102 -176 -83 -172
rect -77 -176 -66 -172
rect -116 -179 -112 -176
rect -175 -185 -128 -181
rect -109 -181 -105 -176
rect -70 -179 -66 -176
rect -109 -185 -82 -181
rect -175 -199 -171 -185
rect -7 -169 9 -165
rect 44 -164 48 -155
rect 31 -168 69 -164
rect 90 -164 94 -155
rect 124 -163 128 -154
rect 282 -114 286 -70
rect 316 -75 320 -70
rect 367 -75 371 -70
rect 413 -75 417 -70
rect 77 -168 116 -164
rect 124 -167 136 -163
rect -21 -184 -16 -179
rect -7 -181 -3 -169
rect 10 -176 16 -172
rect 66 -172 69 -168
rect 124 -171 128 -167
rect 141 -167 142 -163
rect 171 -165 175 -155
rect 21 -176 39 -172
rect 45 -176 63 -172
rect 66 -176 85 -172
rect 91 -176 102 -172
rect 52 -179 56 -176
rect -7 -185 40 -181
rect 59 -181 63 -176
rect 98 -179 102 -176
rect 59 -185 86 -181
rect -183 -245 -179 -239
rect -112 -245 -108 -236
rect -66 -245 -62 -236
rect -52 -245 -47 -191
rect -7 -199 -3 -185
rect 159 -169 175 -165
rect 210 -164 214 -155
rect 197 -168 235 -164
rect 256 -164 260 -155
rect 290 -163 294 -154
rect 447 -114 451 -70
rect 243 -168 282 -164
rect 290 -167 300 -163
rect 145 -184 150 -179
rect 159 -181 163 -169
rect 176 -176 182 -172
rect 232 -172 235 -168
rect 290 -171 294 -167
rect 336 -165 340 -155
rect 187 -176 205 -172
rect 211 -176 229 -172
rect 232 -176 251 -172
rect 257 -176 268 -172
rect 218 -179 222 -176
rect 159 -185 206 -181
rect 225 -181 229 -176
rect 264 -179 268 -176
rect 225 -185 252 -181
rect -15 -245 -11 -239
rect 56 -245 60 -236
rect 102 -245 106 -236
rect 116 -245 121 -191
rect 159 -199 163 -185
rect 324 -169 340 -165
rect 375 -164 379 -155
rect 362 -168 400 -164
rect 421 -164 425 -155
rect 455 -163 459 -154
rect 408 -168 447 -164
rect 455 -167 469 -163
rect 310 -184 315 -179
rect 324 -181 328 -169
rect 341 -176 347 -172
rect 397 -172 400 -168
rect 455 -171 459 -167
rect 352 -176 370 -172
rect 376 -176 394 -172
rect 397 -176 416 -172
rect 422 -176 433 -172
rect 383 -179 387 -176
rect 324 -185 371 -181
rect 390 -181 394 -176
rect 429 -179 433 -176
rect 390 -185 417 -181
rect 151 -245 155 -239
rect 222 -245 226 -236
rect 268 -245 272 -236
rect 282 -245 287 -191
rect 324 -199 328 -185
rect 316 -245 320 -239
rect 387 -245 391 -236
rect 433 -245 437 -236
rect 447 -245 452 -191
rect 497 -245 502 1
rect 525 -211 529 103
rect 558 99 564 100
rect 558 58 564 94
rect 570 99 576 100
rect 570 68 576 94
rect 583 78 589 93
rect 693 77 697 103
rect 752 77 756 103
rect 763 94 822 98
rect 763 77 767 94
rect 818 77 822 94
rect 715 13 718 37
rect 727 28 731 37
rect 775 29 779 37
rect 727 24 774 28
rect 785 11 789 37
rect 826 29 830 37
rect 874 60 877 103
rect 882 11 886 20
rect 720 8 874 11
rect 577 -1 687 3
rect 692 -1 694 3
rect 641 -10 706 -6
rect 694 -14 698 -10
rect 694 -18 724 -14
rect 632 -26 729 -22
rect 564 -34 727 -30
rect 732 -35 742 -31
rect 675 -43 754 -39
rect 732 -52 766 -48
rect 692 -59 778 -55
rect 715 -81 718 -73
rect 727 -75 774 -71
rect 727 -81 731 -75
rect 775 -81 779 -75
rect 785 -81 789 8
rect 882 7 896 11
rect 882 3 886 7
rect 806 -75 830 -71
rect 826 -81 830 -75
rect 693 -112 697 -101
rect 751 -112 755 -101
rect 764 -106 767 -101
rect 818 -106 822 -101
rect 764 -109 822 -106
rect 874 -111 878 -17
rect 925 -111 929 138
rect 1024 127 1028 411
rect 1049 372 1082 376
rect 1137 353 1251 357
rect 1259 299 1263 411
rect 1298 406 1302 412
rect 1362 406 1370 412
rect 1306 357 1310 366
rect 1277 353 1298 357
rect 1306 353 1321 357
rect 1278 291 1283 353
rect 1306 349 1310 353
rect 1213 250 1243 251
rect 1213 246 1247 250
rect 1267 250 1271 259
rect 1252 246 1259 250
rect 1267 246 1286 250
rect 1267 242 1271 246
rect 1259 214 1263 222
rect 1298 214 1302 329
rect 1317 307 1321 353
rect 1414 353 1423 357
rect 1342 318 1346 326
rect 1386 318 1390 326
rect 1342 313 1407 318
rect 1317 303 1341 307
rect 1325 295 1354 299
rect 1324 285 1366 289
rect 1317 275 1379 279
rect 1317 251 1322 275
rect 1342 265 1390 270
rect 1342 261 1346 265
rect 1386 261 1390 265
rect 1374 221 1382 223
rect 1352 214 1356 221
rect 1259 210 1356 214
rect 1376 214 1380 221
rect 1394 214 1398 313
rect 1402 250 1407 313
rect 1431 299 1435 412
rect 1470 406 1474 412
rect 1534 406 1542 412
rect 1478 357 1482 366
rect 1449 353 1470 357
rect 1478 353 1493 357
rect 1450 291 1455 353
rect 1478 349 1482 353
rect 1402 246 1419 250
rect 1439 250 1443 259
rect 1424 246 1431 250
rect 1439 246 1458 250
rect 1439 242 1443 246
rect 1376 210 1398 214
rect 1431 214 1435 222
rect 1470 214 1474 329
rect 1489 307 1493 353
rect 1514 318 1518 326
rect 1558 318 1562 326
rect 1514 313 1576 318
rect 1489 303 1513 307
rect 1497 295 1526 299
rect 1496 285 1538 289
rect 1489 275 1551 279
rect 1489 251 1494 275
rect 1514 265 1562 270
rect 1514 261 1518 265
rect 1558 261 1562 265
rect 1546 221 1554 223
rect 1524 214 1528 221
rect 1431 210 1528 214
rect 1548 214 1552 221
rect 1566 214 1570 313
rect 1548 210 1570 214
rect 1351 203 1356 210
rect 1431 204 1435 210
rect 1594 204 1602 485
rect 1431 203 1602 204
rect 1351 197 1602 203
rect 1060 155 1242 156
rect 1060 147 1402 155
rect 1024 123 1566 127
rect 1024 122 1261 123
rect 873 -112 930 -111
rect 693 -116 930 -112
rect 693 -117 878 -116
rect 544 -166 607 -163
rect 544 -167 617 -166
rect 547 -179 610 -174
rect 616 -179 618 -174
rect 547 -189 608 -184
rect 617 -189 618 -184
rect 626 -194 631 -159
rect 636 -184 641 -159
rect 646 -173 652 -158
rect 547 -199 610 -194
rect 525 -216 786 -211
rect 564 -226 727 -222
rect 632 -238 691 -234
rect 687 -241 691 -238
rect -187 -250 502 -245
rect 447 -400 452 -250
rect 687 -261 691 -246
rect 699 -261 703 -255
rect 711 -261 715 -237
rect 723 -250 727 -226
rect 723 -261 727 -255
rect 760 -261 764 -246
rect 782 -257 786 -216
rect 782 -261 806 -257
rect 788 -267 792 -261
rect 731 -303 736 -299
rect 683 -324 687 -308
rect 683 -350 687 -329
rect 705 -334 709 -308
rect 717 -317 720 -308
rect 757 -317 760 -308
rect 717 -321 760 -317
rect 764 -325 768 -308
rect 764 -343 768 -330
rect 788 -333 792 -307
rect 796 -343 800 -307
rect 764 -347 788 -343
rect 796 -347 811 -343
rect 764 -350 768 -347
rect 731 -363 735 -359
rect 683 -390 687 -370
rect 693 -376 697 -370
rect 705 -400 709 -370
rect 717 -380 721 -370
rect 756 -380 760 -370
rect 717 -384 760 -380
rect 764 -389 768 -370
rect 796 -373 800 -347
rect 788 -400 793 -393
rect 873 -398 877 -117
rect 1024 -180 1028 122
rect 1121 68 1239 69
rect 1121 64 1249 68
rect 1049 7 1069 11
rect 1257 10 1261 122
rect 1296 117 1300 123
rect 1360 117 1368 123
rect 1304 68 1308 77
rect 1275 64 1296 68
rect 1304 64 1319 68
rect 1276 2 1281 64
rect 1304 60 1308 64
rect 1196 -43 1245 -39
rect 1265 -39 1269 -30
rect 1250 -43 1257 -39
rect 1265 -43 1284 -39
rect 1196 -44 1239 -43
rect 1265 -47 1269 -43
rect 1257 -75 1261 -67
rect 1296 -75 1300 40
rect 1315 18 1319 64
rect 1412 64 1421 68
rect 1340 29 1344 37
rect 1384 29 1388 37
rect 1340 24 1405 29
rect 1315 14 1339 18
rect 1323 6 1352 10
rect 1322 -4 1364 0
rect 1315 -14 1377 -10
rect 1315 -38 1320 -14
rect 1340 -24 1388 -19
rect 1340 -28 1344 -24
rect 1384 -28 1388 -24
rect 1372 -68 1380 -66
rect 1350 -75 1354 -68
rect 1257 -79 1354 -75
rect 1374 -75 1378 -68
rect 1392 -75 1396 24
rect 1400 -39 1405 24
rect 1429 10 1433 123
rect 1468 117 1472 123
rect 1532 117 1540 123
rect 1476 68 1480 77
rect 1447 64 1468 68
rect 1476 64 1491 68
rect 1448 2 1453 64
rect 1476 60 1480 64
rect 1400 -43 1417 -39
rect 1437 -39 1441 -30
rect 1422 -43 1429 -39
rect 1437 -43 1456 -39
rect 1437 -47 1441 -43
rect 1374 -79 1396 -75
rect 1429 -75 1433 -67
rect 1468 -75 1472 40
rect 1487 18 1491 64
rect 1512 29 1516 37
rect 1556 29 1560 37
rect 1512 24 1576 29
rect 1487 14 1511 18
rect 1495 6 1524 10
rect 1494 -4 1536 0
rect 1487 -14 1549 -10
rect 1487 -38 1492 -14
rect 1512 -24 1560 -19
rect 1512 -28 1516 -24
rect 1556 -28 1560 -24
rect 1544 -68 1552 -66
rect 1522 -75 1526 -68
rect 1429 -79 1526 -75
rect 1546 -75 1550 -68
rect 1564 -75 1568 24
rect 1546 -79 1568 -75
rect 1349 -86 1354 -79
rect 1429 -85 1433 -79
rect 1594 -85 1602 197
rect 1429 -86 1602 -85
rect 1349 -92 1602 -86
rect 1033 -159 1040 -152
rect 1049 -160 1402 -152
rect 1024 -184 1563 -180
rect 1024 -185 1258 -184
rect 1174 -243 1246 -239
rect 1254 -297 1258 -185
rect 1293 -190 1297 -184
rect 1357 -190 1365 -184
rect 1301 -239 1305 -230
rect 1272 -243 1293 -239
rect 1301 -243 1316 -239
rect 1273 -305 1278 -243
rect 1301 -247 1305 -243
rect 1104 -350 1242 -346
rect 1262 -346 1266 -337
rect 1247 -350 1254 -346
rect 1262 -350 1281 -346
rect 1262 -354 1266 -350
rect 1254 -382 1258 -374
rect 1293 -382 1297 -267
rect 1312 -289 1316 -243
rect 1412 -243 1418 -239
rect 1337 -278 1341 -270
rect 1381 -278 1385 -270
rect 1337 -283 1402 -278
rect 1312 -293 1336 -289
rect 1320 -301 1349 -297
rect 1319 -311 1361 -307
rect 1312 -321 1374 -317
rect 1312 -345 1317 -321
rect 1337 -331 1385 -326
rect 1337 -335 1341 -331
rect 1381 -335 1385 -331
rect 1369 -375 1377 -373
rect 1347 -382 1351 -375
rect 1254 -386 1351 -382
rect 1371 -382 1375 -375
rect 1389 -382 1393 -283
rect 1397 -346 1402 -283
rect 1426 -297 1430 -184
rect 1465 -190 1469 -184
rect 1529 -190 1537 -184
rect 1473 -239 1477 -230
rect 1444 -243 1465 -239
rect 1473 -243 1488 -239
rect 1445 -305 1450 -243
rect 1473 -247 1477 -243
rect 1397 -350 1414 -346
rect 1434 -346 1438 -337
rect 1419 -350 1426 -346
rect 1434 -350 1453 -346
rect 1434 -354 1438 -350
rect 1371 -386 1393 -382
rect 1426 -382 1430 -374
rect 1465 -382 1469 -267
rect 1484 -289 1488 -243
rect 1509 -278 1513 -270
rect 1553 -278 1557 -270
rect 1509 -283 1573 -278
rect 1484 -293 1508 -289
rect 1492 -301 1521 -297
rect 1491 -311 1533 -307
rect 1484 -321 1546 -317
rect 1484 -345 1489 -321
rect 1509 -331 1557 -326
rect 1509 -335 1513 -331
rect 1553 -335 1557 -331
rect 1541 -375 1549 -373
rect 1519 -382 1523 -375
rect 1426 -386 1523 -382
rect 1543 -382 1547 -375
rect 1561 -382 1565 -283
rect 1543 -386 1565 -382
rect 1346 -393 1351 -386
rect 1426 -393 1430 -386
rect 1593 -393 1602 -92
rect 872 -400 877 -398
rect 447 -404 877 -400
rect 872 -555 877 -404
rect 1345 -399 1602 -393
rect 1097 -541 1102 -439
rect 1114 -529 1119 -441
rect 1130 -515 1135 -441
rect 1149 -499 1154 -442
rect 1168 -478 1173 -441
rect 1189 -468 1194 -441
rect 1205 -457 1210 -439
rect 1345 -555 1351 -399
rect 1430 -400 1602 -399
rect 872 -560 1351 -555
<< m2contact >>
rect 795 865 802 871
rect 867 881 872 887
rect 878 881 884 887
rect 867 862 872 868
rect 878 840 884 849
rect 795 828 802 834
rect 723 813 729 822
rect 595 797 600 802
rect 681 794 691 802
rect 657 785 662 790
rect 646 768 651 773
rect 711 768 717 773
rect 583 758 588 763
rect 735 758 741 764
rect 569 749 574 754
rect 698 749 704 754
rect 636 741 641 746
rect 747 741 752 746
rect 711 732 717 737
rect 735 723 741 729
rect 747 714 752 719
rect 626 705 631 710
rect 808 705 813 710
rect 558 696 563 701
rect 820 696 826 701
rect 667 687 673 692
rect 820 678 826 683
rect 698 669 704 674
rect 808 660 813 665
rect 681 650 691 658
rect 723 576 729 585
rect 794 638 801 646
rect 794 583 802 591
rect 878 625 883 632
rect 867 596 873 603
rect 867 571 873 578
rect 878 572 883 577
rect 773 421 779 426
rect 797 421 803 426
rect 858 422 864 427
rect 713 370 719 376
rect 945 372 950 377
rect 583 360 589 365
rect 686 359 692 365
rect 646 351 652 356
rect 636 335 642 340
rect 701 334 706 340
rect 570 324 576 329
rect 725 324 731 330
rect 558 316 564 321
rect 737 317 742 322
rect 626 309 632 314
rect 749 308 755 314
rect 701 299 706 306
rect 725 289 731 296
rect 738 278 743 283
rect 667 268 676 273
rect 749 257 755 263
rect 686 248 692 254
rect 713 227 718 232
rect 773 204 778 209
rect 799 205 804 210
rect 858 205 863 210
rect -141 83 -136 88
rect -95 83 -90 88
rect -33 84 -27 90
rect -151 75 -146 80
rect 27 83 32 88
rect 73 83 78 88
rect 17 75 22 80
rect 137 83 142 88
rect -132 55 -127 60
rect -86 55 -81 60
rect 193 83 198 88
rect 239 83 244 88
rect 183 75 188 80
rect 301 83 306 89
rect 36 55 41 60
rect 82 55 87 60
rect 358 83 363 88
rect 404 83 409 88
rect 1080 722 1089 733
rect 1409 723 1420 732
rect 1221 640 1229 646
rect 1256 640 1261 646
rect 1277 641 1282 646
rect 1283 572 1289 579
rect 1148 533 1154 538
rect 1252 534 1257 539
rect 1291 533 1297 539
rect 1409 639 1419 646
rect 1428 640 1433 646
rect 1324 582 1330 588
rect 1323 571 1329 578
rect 1321 534 1327 539
rect 1449 641 1454 646
rect 1455 572 1461 579
rect 1424 534 1429 539
rect 1463 533 1469 539
rect 1496 582 1502 588
rect 1495 571 1501 578
rect 1493 534 1499 539
rect 1067 435 1078 445
rect 1404 435 1415 444
rect 348 75 353 80
rect 470 83 476 89
rect 202 55 207 60
rect 248 55 253 60
rect 367 55 372 60
rect 413 55 418 60
rect -142 -168 -137 -163
rect -96 -168 -91 -163
rect -34 -167 -28 -161
rect -152 -176 -147 -171
rect 26 -168 31 -163
rect 72 -168 77 -163
rect 16 -176 21 -171
rect 136 -168 141 -163
rect -133 -196 -128 -191
rect -87 -196 -82 -191
rect 192 -168 197 -163
rect 238 -168 243 -163
rect 182 -176 187 -171
rect 300 -168 305 -162
rect 35 -196 40 -191
rect 81 -196 86 -191
rect 357 -168 362 -163
rect 403 -168 408 -163
rect 347 -176 352 -171
rect 469 -168 475 -162
rect 201 -196 206 -191
rect 247 -196 252 -191
rect 366 -196 371 -191
rect 412 -196 417 -191
rect 557 94 564 99
rect 570 94 577 99
rect 583 93 590 98
rect 583 72 590 78
rect 570 62 577 68
rect 558 52 565 58
rect 774 24 779 29
rect 714 8 720 13
rect 826 24 831 29
rect 569 -2 577 3
rect 687 -2 692 4
rect 635 -11 641 -5
rect 626 -26 632 -20
rect 558 -35 564 -29
rect 727 -35 732 -30
rect 667 -43 675 -38
rect 727 -52 732 -47
rect 686 -59 692 -54
rect 714 -73 719 -68
rect 774 -75 780 -70
rect 896 7 902 12
rect 799 -75 806 -70
rect 1044 371 1049 377
rect 1082 371 1089 377
rect 1129 350 1137 357
rect 1251 352 1256 358
rect 1272 353 1277 358
rect 1278 284 1284 291
rect 1201 243 1213 252
rect 1247 246 1252 251
rect 1286 245 1292 251
rect 1404 351 1414 358
rect 1423 352 1428 358
rect 1319 294 1325 300
rect 1318 283 1324 290
rect 1316 246 1322 251
rect 1444 353 1449 358
rect 1450 284 1456 291
rect 1419 246 1424 251
rect 1458 245 1464 251
rect 1491 294 1497 300
rect 1490 283 1496 290
rect 1488 246 1494 251
rect 1045 140 1060 160
rect 1402 146 1413 155
rect 625 -159 631 -154
rect 635 -159 642 -154
rect 646 -158 652 -152
rect 538 -168 544 -161
rect 607 -166 617 -161
rect 538 -179 547 -174
rect 610 -179 616 -172
rect 538 -189 547 -184
rect 608 -189 617 -184
rect 645 -180 653 -173
rect 634 -190 641 -184
rect 538 -199 547 -194
rect 610 -199 619 -194
rect 625 -200 631 -194
rect 557 -227 564 -222
rect 624 -239 632 -234
rect 710 -237 716 -232
rect 686 -246 691 -241
rect 699 -255 704 -250
rect 759 -246 764 -241
rect 722 -255 727 -250
rect 736 -303 742 -298
rect 681 -329 687 -324
rect 704 -339 709 -334
rect 764 -330 770 -325
rect 787 -339 792 -333
rect 811 -347 816 -342
rect 735 -364 740 -357
rect 683 -396 688 -390
rect 763 -396 770 -389
rect 1112 63 1121 69
rect 1249 63 1254 69
rect 1037 4 1049 12
rect 1069 6 1075 12
rect 1270 64 1275 69
rect 1276 -5 1282 2
rect 1186 -45 1196 -38
rect 1245 -43 1250 -38
rect 1284 -44 1290 -38
rect 1402 62 1412 69
rect 1421 63 1426 69
rect 1317 5 1323 11
rect 1316 -6 1322 1
rect 1314 -43 1320 -38
rect 1442 64 1447 69
rect 1448 -5 1454 2
rect 1417 -43 1422 -38
rect 1456 -44 1462 -38
rect 1489 5 1495 11
rect 1488 -6 1494 1
rect 1486 -43 1492 -38
rect 1040 -162 1049 -150
rect 1402 -161 1413 -152
rect 1166 -245 1174 -237
rect 1246 -244 1251 -238
rect 1267 -243 1272 -238
rect 1273 -312 1279 -305
rect 1096 -352 1104 -345
rect 1242 -350 1247 -345
rect 1281 -351 1287 -345
rect 1402 -245 1412 -238
rect 1418 -244 1423 -238
rect 1314 -302 1320 -296
rect 1313 -313 1319 -306
rect 1311 -350 1317 -345
rect 1439 -243 1444 -238
rect 1445 -312 1451 -305
rect 1414 -350 1419 -345
rect 1453 -351 1459 -345
rect 1486 -302 1492 -296
rect 1485 -313 1491 -306
rect 1483 -350 1489 -345
rect 1097 -439 1102 -433
rect 1114 -441 1119 -435
rect 1130 -441 1135 -435
rect 1149 -442 1154 -436
rect 1167 -441 1174 -436
rect 1188 -441 1195 -431
rect 1204 -439 1210 -431
rect 1203 -465 1210 -457
rect 1189 -476 1196 -468
rect 1168 -486 1175 -478
rect 1148 -507 1155 -499
rect 1129 -523 1136 -515
rect 1112 -537 1119 -529
rect 1096 -549 1103 -541
<< metal2 >>
rect 867 868 872 881
rect 796 834 801 865
rect 878 849 882 881
rect 558 701 564 812
rect 570 754 576 812
rect 574 749 576 754
rect 563 696 564 701
rect 558 321 564 696
rect -228 195 353 199
rect -228 -51 -223 195
rect -151 80 -146 195
rect -151 74 -146 75
rect -141 60 -136 83
rect -95 60 -90 83
rect -141 55 -132 60
rect -95 55 -86 60
rect -32 -23 -28 84
rect 17 80 22 195
rect 27 60 32 83
rect 73 60 78 83
rect 27 55 36 60
rect 73 55 82 60
rect 137 -13 141 83
rect 183 80 188 195
rect 193 60 198 83
rect 239 60 244 83
rect 193 55 202 60
rect 239 55 248 60
rect 301 -4 305 83
rect 348 80 353 195
rect 558 99 564 316
rect 570 329 576 749
rect 570 99 576 324
rect 583 763 589 812
rect 588 758 589 763
rect 583 365 589 758
rect 583 98 589 360
rect 595 802 600 812
rect 358 60 363 83
rect 595 88 600 797
rect 476 84 600 88
rect 404 60 409 83
rect 473 72 583 77
rect 358 55 367 60
rect 404 55 413 60
rect 473 -4 478 72
rect 301 -8 478 -4
rect 487 62 570 67
rect 487 -13 491 62
rect 137 -17 491 -13
rect 497 52 558 57
rect 497 -23 501 52
rect -32 -28 501 -23
rect 558 -29 564 52
rect 570 3 576 62
rect -228 -56 351 -51
rect -152 -171 -148 -56
rect -142 -191 -137 -168
rect -96 -191 -91 -168
rect -142 -196 -133 -191
rect -96 -196 -87 -191
rect -33 -274 -29 -167
rect 16 -171 20 -56
rect 26 -191 31 -168
rect 72 -191 77 -168
rect 26 -196 35 -191
rect 72 -196 81 -191
rect 136 -264 140 -168
rect 182 -171 186 -56
rect 346 -57 351 -56
rect 192 -191 197 -168
rect 238 -191 243 -168
rect 192 -196 201 -191
rect 238 -196 247 -191
rect 300 -255 304 -168
rect 347 -171 351 -57
rect 357 -191 362 -168
rect 475 -167 538 -163
rect 403 -191 408 -168
rect 472 -179 538 -174
rect 357 -196 366 -191
rect 403 -196 412 -191
rect 472 -255 477 -179
rect 300 -259 477 -255
rect 486 -189 538 -184
rect 486 -264 490 -189
rect 136 -268 490 -264
rect 496 -199 538 -194
rect 496 -274 500 -199
rect 558 -222 564 -35
rect -33 -279 500 -274
rect 558 -542 564 -227
rect 570 -530 576 -2
rect 583 -515 589 72
rect 595 -502 600 84
rect 626 710 631 812
rect 626 314 631 705
rect 636 746 641 812
rect 636 340 641 741
rect 646 773 652 812
rect 651 768 652 773
rect 646 356 652 768
rect 626 -20 631 309
rect 636 -5 641 335
rect 626 -154 631 -26
rect 636 -154 641 -11
rect 646 -152 652 351
rect 657 790 662 812
rect 657 -163 662 785
rect 667 273 673 687
rect 682 658 690 794
rect 698 674 704 749
rect 711 737 717 768
rect 724 585 728 813
rect 735 729 741 758
rect 747 719 752 741
rect 808 665 812 705
rect 820 683 825 696
rect 795 591 800 638
rect 868 578 872 596
rect 724 571 728 576
rect 878 577 882 625
rect 878 571 882 572
rect 779 422 797 426
rect 803 422 858 426
rect 714 376 718 377
rect 950 372 1044 376
rect 667 -38 675 268
rect 686 254 692 359
rect 701 306 705 334
rect 714 232 718 370
rect 726 296 730 324
rect 742 317 743 321
rect 737 283 743 317
rect 737 278 738 283
rect 750 263 754 308
rect 1053 250 1057 758
rect 1070 445 1074 758
rect 1083 733 1087 758
rect 1048 238 1061 250
rect 778 205 799 209
rect 804 205 858 209
rect 1053 160 1057 238
rect 779 24 826 28
rect 667 -153 675 -43
rect 687 -54 691 -2
rect 715 -68 718 8
rect 902 7 1037 11
rect 727 -47 731 -35
rect 780 -75 799 -71
rect 806 -75 807 -71
rect 666 -161 1040 -153
rect 617 -166 662 -163
rect 607 -167 662 -166
rect 608 -179 610 -174
rect 616 -179 645 -174
rect 617 -189 634 -184
rect 608 -199 610 -194
rect 619 -199 625 -194
rect 626 -234 631 -200
rect 626 -481 631 -239
rect 636 -469 641 -190
rect 646 -459 652 -180
rect 657 -447 662 -167
rect 667 -202 675 -161
rect 667 -206 715 -202
rect 711 -232 715 -206
rect 691 -246 759 -242
rect 704 -255 722 -251
rect 736 -326 741 -303
rect 687 -329 764 -326
rect 709 -339 787 -334
rect 1053 -343 1057 140
rect 1070 12 1074 435
rect 1083 377 1087 722
rect 816 -347 1057 -343
rect 1097 -345 1102 758
rect 1114 162 1119 758
rect 1130 357 1135 758
rect 1149 538 1154 758
rect 1113 157 1120 162
rect 1114 69 1119 157
rect 735 -391 739 -364
rect 688 -395 763 -391
rect 1097 -433 1102 -352
rect 1114 -435 1119 63
rect 1130 -435 1135 350
rect 1149 -436 1154 533
rect 1168 -237 1173 758
rect 1189 55 1194 758
rect 1205 252 1210 758
rect 1223 646 1228 758
rect 1411 646 1418 723
rect 1261 641 1277 645
rect 1188 49 1196 55
rect 1189 -38 1194 49
rect 1168 -436 1173 -245
rect 1189 -431 1194 -45
rect 1205 -431 1210 243
rect 1223 -447 1228 640
rect 1433 641 1449 645
rect 1253 583 1324 587
rect 1253 539 1257 583
rect 1425 583 1496 587
rect 1289 573 1323 577
rect 1425 539 1429 583
rect 1461 573 1495 577
rect 1297 534 1321 538
rect 1469 534 1493 538
rect 1406 358 1413 435
rect 1256 353 1272 357
rect 1428 353 1444 357
rect 1248 295 1319 299
rect 1248 251 1252 295
rect 1420 295 1491 299
rect 1284 285 1318 289
rect 1420 251 1424 295
rect 1456 285 1490 289
rect 1292 246 1316 250
rect 1464 246 1488 250
rect 1404 69 1411 146
rect 1254 64 1270 68
rect 1426 64 1442 68
rect 1246 6 1317 10
rect 1246 -38 1250 6
rect 1418 6 1489 10
rect 1282 -4 1316 0
rect 1418 -38 1422 6
rect 1454 -4 1488 0
rect 1290 -43 1314 -39
rect 1462 -43 1486 -39
rect 1404 -238 1411 -161
rect 1251 -243 1267 -239
rect 1423 -243 1439 -239
rect 1243 -301 1314 -297
rect 1243 -345 1247 -301
rect 1415 -301 1486 -297
rect 1279 -311 1313 -307
rect 1415 -345 1419 -301
rect 1451 -311 1485 -307
rect 1287 -350 1311 -346
rect 1459 -350 1483 -346
rect 657 -452 1228 -447
rect 646 -464 1203 -459
rect 636 -474 1189 -469
rect 626 -486 1168 -481
rect 595 -507 1148 -502
rect 583 -522 1129 -515
rect 570 -535 1112 -530
rect 558 -547 1096 -542
<< labels >>
rlabel metal1 -154 77 -154 77 1 clk
rlabel metal1 -174 2 -174 2 1 gnd
rlabel metal1 -81 187 -81 187 5 vdd
rlabel metal1 -127 187 -127 187 5 vdd
rlabel metal1 -170 188 -170 188 5 vdd
rlabel metal1 -187 68 -185 71 3 a0_in
rlabel metal1 -36 85 -33 87 1 a0
rlabel metal1 14 77 14 77 1 clk
rlabel metal1 -6 2 -6 2 1 gnd
rlabel metal1 87 187 87 187 5 vdd
rlabel metal1 41 187 41 187 5 vdd
rlabel metal1 -2 188 -2 188 5 vdd
rlabel metal1 -20 67 -14 72 1 a1_in
rlabel metal1 132 84 136 88 1 a1
rlabel metal1 180 77 180 77 1 clk
rlabel metal1 160 2 160 2 1 gnd
rlabel metal1 253 187 253 187 5 vdd
rlabel metal1 207 187 207 187 5 vdd
rlabel metal1 164 188 164 188 5 vdd
rlabel space 146 67 152 73 1 a2_in
rlabel space 298 83 303 89 1 a2
rlabel metal1 345 77 345 77 1 clk
rlabel metal1 325 2 325 2 1 gnd
rlabel metal1 418 187 418 187 5 vdd
rlabel metal1 372 187 372 187 5 vdd
rlabel metal1 329 188 329 188 5 vdd
rlabel metal1 311 67 316 72 1 a3_in
rlabel metal1 463 84 467 88 1 a3
rlabel metal2 503 84 508 88 1 a3
rlabel metal2 504 73 508 77 1 a2
rlabel space 504 61 509 67 1 a1
rlabel metal1 -155 -174 -155 -174 1 clk
rlabel metal1 -175 -249 -175 -249 1 gnd
rlabel metal1 -82 -64 -82 -64 5 vdd
rlabel metal1 -128 -64 -128 -64 5 vdd
rlabel metal1 -171 -63 -171 -63 5 vdd
rlabel metal1 13 -174 13 -174 1 clk
rlabel metal1 -7 -249 -7 -249 1 gnd
rlabel metal1 86 -64 86 -64 5 vdd
rlabel metal1 40 -64 40 -64 5 vdd
rlabel metal1 -3 -63 -3 -63 5 vdd
rlabel metal1 179 -174 179 -174 1 clk
rlabel metal1 159 -249 159 -249 1 gnd
rlabel metal1 252 -64 252 -64 5 vdd
rlabel metal1 206 -64 206 -64 5 vdd
rlabel metal1 163 -63 163 -63 5 vdd
rlabel metal1 344 -174 344 -174 1 clk
rlabel metal1 324 -249 324 -249 1 gnd
rlabel metal1 417 -64 417 -64 5 vdd
rlabel metal1 371 -64 371 -64 5 vdd
rlabel metal1 328 -63 328 -63 5 vdd
rlabel metal1 -189 -184 -182 -179 3 b0_in
rlabel space -38 -168 -34 -163 1 b0
rlabel metal1 -21 -184 -15 -179 1 b1_in
rlabel space 131 -168 135 -162 1 b1
rlabel metal1 145 -184 150 -179 1 b2_in
rlabel metal1 296 -167 299 -163 1 b2
rlabel metal1 310 -184 315 -179 1 b3_in
rlabel metal1 462 -167 466 -163 1 b3
rlabel metal2 498 -167 503 -163 1 b3
rlabel metal2 498 -178 503 -174 1 b2
rlabel metal2 498 -189 503 -185 1 b1
rlabel metal2 501 -199 506 -195 1 b0
rlabel metal1 668 -26 674 -22 1 b0
rlabel metal1 668 -1 672 3 1 a1
rlabel metal1 681 360 686 364 1 a2
rlabel metal1 682 351 687 355 1 b2
rlabel metal1 683 335 687 339 1 b1
rlabel metal1 683 325 687 329 1 a1
rlabel metal1 685 309 689 313 1 b0
rlabel metal1 685 268 690 273 1 cin
rlabel metal1 942 372 949 376 7 c3
rlabel metal1 930 141 930 141 1 gnd
rlabel metal1 670 797 675 802 1 a3
rlabel metal1 670 768 676 773 1 b2
rlabel metal1 670 759 676 764 1 a2
rlabel metal1 670 741 676 746 1 b1
rlabel metal1 666 785 671 790 1 b3
rlabel metal1 666 749 671 754 1 a1
rlabel metal1 675 706 680 710 1 b0
rlabel metal1 676 696 681 700 1 a0
rlabel metal1 675 687 681 692 1 cin
rlabel metal1 1007 817 1012 821 1 cout
rlabel metal1 956 942 963 945 5 vdd
rlabel space 521 52 526 58 1 a0
rlabel metal1 689 -259 689 -259 1 b0
rlabel metal1 702 -259 702 -259 1 a0
rlabel metal1 713 -259 713 -259 1 cin
rlabel metal1 725 -259 725 -259 1 a0
rlabel metal1 763 -259 763 -259 1 b0
rlabel metal1 793 -259 793 -259 5 vdd
rlabel metal1 684 -331 684 -331 1 n010
rlabel metal2 741 -328 741 -328 1 n010
rlabel metal1 793 -402 793 -402 1 gnd
rlabel metal2 738 -393 738 -393 1 n010
rlabel metal1 777 -345 777 -345 1 n010
rlabel metal1 809 -345 809 -345 1 c1
rlabel metal1 707 -381 707 -381 1 gnd
rlabel metal1 860 -116 867 -113 1 gnd
rlabel metal1 686 0 689 3 3 a1
rlabel metal1 687 -10 691 -6 3 b1
rlabel metal1 688 -26 691 -22 3 b0
rlabel metal1 688 -43 691 -39 3 cin
rlabel m2contact 669 -43 674 -39 1 cin
rlabel metal1 890 7 895 11 1 c2
rlabel metal1 852 103 861 107 5 vdd
rlabel metal1 915 516 915 516 5 vdd
rlabel metal1 1259 -384 1259 -384 1 gnd
rlabel metal1 1259 -182 1259 -182 5 vdd
rlabel metal1 1300 -384 1300 -384 1 gnd
rlabel metal1 1298 -181 1298 -181 5 vdd
rlabel metal1 1431 -384 1431 -384 1 gnd
rlabel metal1 1431 -182 1431 -182 5 vdd
rlabel metal1 1472 -384 1472 -384 1 gnd
rlabel metal1 1470 -181 1470 -181 5 vdd
rlabel metal1 1564 -283 1573 -278 1 s0_out
rlabel metal1 1262 -77 1262 -77 1 gnd
rlabel metal1 1262 125 1262 125 5 vdd
rlabel metal1 1303 -77 1303 -77 1 gnd
rlabel metal1 1301 126 1301 126 5 vdd
rlabel metal1 1434 -77 1434 -77 1 gnd
rlabel metal1 1434 125 1434 125 5 vdd
rlabel metal1 1475 -77 1475 -77 1 gnd
rlabel metal1 1473 126 1473 126 5 vdd
rlabel space 1568 23 1576 30 7 s1_out
rlabel metal1 1264 212 1264 212 1 gnd
rlabel metal1 1264 414 1264 414 5 vdd
rlabel metal1 1305 212 1305 212 1 gnd
rlabel metal1 1303 415 1303 415 5 vdd
rlabel metal1 1436 212 1436 212 1 gnd
rlabel metal1 1436 414 1436 414 5 vdd
rlabel metal1 1477 212 1477 212 1 gnd
rlabel metal1 1475 415 1475 415 5 vdd
rlabel metal1 1568 313 1573 318 1 s2_out
rlabel metal1 1269 500 1269 500 1 gnd
rlabel metal1 1269 702 1269 702 5 vdd
rlabel metal1 1310 500 1310 500 1 gnd
rlabel metal1 1308 703 1308 703 5 vdd
rlabel metal1 1441 500 1441 500 1 gnd
rlabel metal1 1441 702 1441 702 5 vdd
rlabel metal1 1482 500 1482 500 1 gnd
rlabel metal1 1480 703 1480 703 5 vdd
rlabel space 1572 600 1579 607 1 s3_out
<< end >>
