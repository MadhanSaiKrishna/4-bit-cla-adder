magic
tech scmos
timestamp 1733158314
<< nwell >>
rect 0 -1 66 52
rect 72 -1 98 52
rect 105 0 129 52
<< ntransistor >>
rect 11 -57 13 -37
rect 23 -57 25 -37
rect 35 -57 37 -37
rect 47 -57 49 -37
rect 84 -57 86 -37
rect 116 -80 118 -60
<< ptransistor >>
rect 11 5 13 45
rect 23 5 25 45
rect 35 5 37 45
rect 47 5 49 45
rect 84 5 86 45
rect 116 6 118 46
<< ndiffusion >>
rect 10 -57 11 -37
rect 13 -57 14 -37
rect 22 -57 23 -37
rect 25 -57 26 -37
rect 34 -57 35 -37
rect 37 -57 38 -37
rect 46 -57 47 -37
rect 49 -57 50 -37
rect 83 -57 84 -37
rect 86 -57 87 -37
rect 115 -80 116 -60
rect 118 -80 119 -60
<< pdiffusion >>
rect 10 5 11 45
rect 13 5 14 45
rect 22 5 23 45
rect 25 5 26 45
rect 34 5 35 45
rect 37 5 38 45
rect 46 5 47 45
rect 49 5 50 45
rect 83 5 84 45
rect 86 5 87 45
rect 115 6 116 46
rect 118 6 119 46
<< ndcontact >>
rect 6 -57 10 -37
rect 14 -57 22 -37
rect 26 -57 34 -37
rect 38 -57 46 -37
rect 50 -57 54 -37
rect 79 -57 83 -37
rect 87 -57 91 -37
rect 111 -80 115 -60
rect 119 -80 123 -60
<< pdcontact >>
rect 6 5 10 45
rect 14 5 22 45
rect 26 5 34 45
rect 38 5 46 45
rect 50 5 54 45
rect 79 5 83 45
rect 87 5 91 45
rect 111 6 115 46
rect 119 6 123 46
<< polysilicon >>
rect 11 45 13 48
rect 23 45 25 48
rect 35 45 37 48
rect 47 45 49 48
rect 84 45 86 48
rect 116 46 118 52
rect 11 -37 13 5
rect 23 -37 25 5
rect 35 -37 37 5
rect 47 -37 49 5
rect 84 -37 86 5
rect 11 -62 13 -57
rect 23 -62 25 -57
rect 35 -61 37 -57
rect 47 -61 49 -57
rect 84 -61 86 -57
rect 116 -60 118 6
rect 116 -84 118 -80
<< polycontact >>
rect 10 48 14 52
rect 22 48 26 52
rect 34 48 38 52
rect 46 48 50 52
rect 83 48 87 52
rect 111 -34 116 -30
<< metal1 >>
rect 10 72 14 79
rect 10 52 14 67
rect 22 52 26 58
rect 34 52 38 79
rect 46 63 50 79
rect 46 52 50 58
rect 83 52 87 67
rect 105 52 129 56
rect 111 46 115 52
rect 54 10 59 14
rect 6 -11 10 5
rect 6 -37 10 -16
rect 28 -21 32 5
rect 40 -4 43 5
rect 80 -4 83 5
rect 40 -8 83 -4
rect 87 -12 91 5
rect 87 -30 91 -17
rect 111 -20 115 6
rect 119 -30 123 6
rect 87 -34 111 -30
rect 119 -34 139 -30
rect 87 -37 91 -34
rect 54 -50 58 -46
rect 6 -77 10 -57
rect 16 -63 20 -57
rect 28 -87 32 -57
rect 40 -67 44 -57
rect 79 -67 83 -57
rect 40 -71 83 -67
rect 87 -76 91 -57
rect 119 -60 123 -34
rect 111 -87 116 -80
rect 5 -91 129 -87
<< m2contact >>
rect 9 67 14 72
rect 22 58 27 63
rect 82 67 87 72
rect 45 58 50 63
rect 59 10 65 15
rect 4 -16 10 -11
rect 27 -26 32 -21
rect 87 -17 93 -12
rect 110 -26 115 -20
rect 58 -51 63 -44
rect 6 -83 11 -77
rect 86 -83 93 -76
<< metal2 >>
rect 14 67 82 71
rect 27 58 45 62
rect 59 -13 64 10
rect 10 -16 87 -13
rect 32 -26 110 -21
rect 58 -78 62 -51
rect 11 -82 86 -78
<< labels >>
rlabel metal1 12 54 12 54 1 b0
rlabel metal1 25 54 25 54 1 a0
rlabel metal1 36 54 36 54 1 cin
rlabel metal1 48 54 48 54 1 a0
rlabel metal1 86 54 86 54 1 b0
rlabel metal1 116 54 116 54 5 vdd
rlabel metal1 7 -18 7 -18 1 n010
rlabel metal2 64 -15 64 -15 1 n010
rlabel metal1 116 -89 116 -89 1 gnd
rlabel metal2 61 -80 61 -80 1 n010
rlabel metal1 100 -32 100 -32 1 n010
rlabel metal1 132 -32 132 -32 1 c1
rlabel metal1 30 -68 30 -68 1 gnd
<< end >>
