* SPICE3 file created from carry_one.ext - technology: scmos
.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY = 1.8
.param LAMBDA=0.09u
.global gnd vdd
Vdd vdd gnd 'SUPPLY'

V1 A0_in gnd pulse 0 1.8 0u 10p 10p 0.1u 0.3u
V2 B0_in gnd pulse 0 1.8 0.3u 10p 10p 0.1u 0.3u
V3 A1_in gnd pulse 0 1.8 0.5u 10p 10p 0.01u 0.03u
V4 B1_in gnd pulse 0 1.8 0u 10p 10p 0.02u 0.03u
V5 A2_in gnd pulse 0 1.8 0.5u 10p 10p 0.1u 0.3u
V6 B2_in gnd pulse 0 1.8 0u 10p 10p 0.1u 0.3u
V7 A3_in gnd pulse 0 1.8 0.5u 10p 10p 0.01u 0.03u
V8 B3_in gnd pulse 0 1.8 0u 10p 10p 0.02u 0.07u

V9 clk gnd pulse 0 1.8 0.03u 10p 10p 60n 100n


V10 Cin gnd dc 0


M1000 a_n7_12# a1_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=7200 ps=3200
M1001 gnd clk a_374_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1002 a_718_n123# a_716_n126# a_706_n123# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=200 ps=60
M1003 a_759_164# a0 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1004 a_723_455# b2 a_711_164# w_686_449# CMOSP w=40 l=2
+  ad=1000 pd=290 as=600 ps=190
M1005 a_817_889# b0 a_853_889# w_902_883# CMOSP w=40 l=2
+  ad=1000 pd=290 as=600 ps=190
M1006 a_n125_n236# a_n176_n239# a_n132_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1007 n010 a0 a_714_n308# w_677_n314# CMOSP w=40 l=2
+  ad=600 pd=270 as=600 ps=190
M1008 a_699_164# a2 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1009 a1 a_83_15# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1010 a_742_n123# b0 a_730_n123# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=500 ps=170
M1011 a_721_551# a3 a_733_889# w_941_883# CMOSP w=40 l=2
+  ad=600 pd=190 as=1000 ps=290
M1012 c2 a_718_50# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1013 a_159_96# a_151_67# vdd w_145_88# CMOSP w=80 l=2
+  ad=800 pd=180 as=14800 ps=6020
M1014 a_255_n236# clk a_248_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1015 a_159_12# a_151_67# gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1016 a_37_15# clk vdd w_29_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1017 a_706_50# a1 vdd w_693_44# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1018 vdd a0 a_829_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1019 a_n85_15# a_n131_15# vdd w_n93_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1020 gnd a_n131_15# a_n78_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1021 a_209_n236# a_158_n239# a_202_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1022 a_82_n236# a_36_n236# vdd w_74_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1023 a_n86_n236# a_n132_n236# vdd w_n94_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1024 cout a_721_551# vdd w_985_824# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1025 a_730_n123# b1 a_718_n123# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 a_83_15# a_37_15# vdd w_75_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1027 a_781_889# b1 a_769_889# w_692_883# CMOSP w=40 l=2
+  ad=1000 pd=290 as=400 ps=100
M1028 a3 a_414_15# vdd w_438_91# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1029 a_771_164# b0 a_759_164# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=0 ps=0
M1030 a_735_455# b1 a_723_455# w_686_449# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1031 a_159_12# clk a_159_96# w_145_88# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1032 a_723_455# b1 a_771_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=1000 ps=290
M1033 a_44_15# a_n7_12# a_37_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1034 a_n8_n155# b1_in vdd w_n22_n163# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1035 a_733_551# b3 a_721_551# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=300 ps=110
M1036 gnd a_37_15# a_90_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1037 a_754_n123# a0 a_742_n123# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1038 a_718_50# b1 a_706_50# w_693_44# CMOSP w=40 l=2
+  ad=600 pd=190 as=0 ps=0
M1039 c3 a_711_164# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1040 a_n78_15# clk a_n85_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1041 a_367_n236# clk vdd w_359_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1042 b1 a_82_n236# vdd w_106_n160# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1043 a_n8_n239# clk a_n8_n155# w_n22_n163# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1044 a_203_15# clk vdd w_195_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1045 b1 a_82_n236# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1046 a_249_15# a_203_15# vdd w_241_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1047 a_90_15# clk a_83_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1048 a_368_15# clk vdd w_360_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1049 a0 a_n85_15# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1050 gnd a_202_n236# a_255_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 a_771_164# b0 a_807_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=300 ps=110
M1052 gnd clk a_209_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 a2 a_249_15# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1054 gnd clk a_44_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 gnd a_367_n236# a_420_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1056 a_730_50# b1 a_718_50# w_693_44# CMOSP w=40 l=2
+  ad=1000 pd=290 as=0 ps=0
M1057 a_711_164# a2 a_723_164# Gnd CMOSN w=20 l=2
+  ad=300 pd=110 as=500 ps=170
M1058 a_690_n370# b0 n010 Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=300 ps=150
M1059 a_807_455# a0 a_771_455# w_686_449# CMOSP w=40 l=2
+  ad=600 pd=190 as=0 ps=0
M1060 a_210_15# a_159_12# a_203_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1061 a_256_15# clk a_249_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1062 a_781_551# a2 a_733_551# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=0 ps=0
M1063 a_n175_12# clk a_n175_96# w_n189_88# CMOSP w=80 l=2
+  ad=400 pd=170 as=800 ps=180
M1064 a_324_96# a3_in vdd w_310_88# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1065 a_375_15# a_324_12# a_368_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1066 a_853_551# cin gnd Gnd CMOSN w=20 l=2
+  ad=300 pd=110 as=0 ps=0
M1067 a_158_n239# b2_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1068 a_766_n123# cin a_754_n123# Gnd CMOSN w=20 l=2
+  ad=300 pd=110 as=0 ps=0
M1069 a_742_50# b0 a_730_50# w_693_44# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1070 a_324_12# a3_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1071 vdd a1 a_735_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 a_771_455# a1 a_723_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 a_420_n236# clk a_413_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1074 gnd clk a_210_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 a_733_889# b3 a_721_551# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 a_745_551# b2 a_733_551# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1077 a_733_551# b2 a_781_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 a_323_n239# b3_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1079 a_n132_n236# clk vdd w_n140_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1080 a_723_164# b2 a_711_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 gnd a_203_15# a_256_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 a_n175_96# a0_in vdd w_n189_88# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 a_324_12# clk a_324_96# w_310_88# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1084 gnd clk a_375_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 a_690_n308# b0 n010 w_677_n314# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1086 vdd a0 a_742_50# w_693_44# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 a_n175_12# a0_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1088 a_43_n236# a_n8_n239# a_36_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1089 a_248_n236# a_202_n236# vdd w_240_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1090 vdd cin a_807_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 a_202_n236# clk vdd w_194_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1092 a_730_n123# a0 a_766_n123# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 c2 a_718_50# vdd w_870_16# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1094 a_781_889# a2 a_733_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 a_817_551# b1 a_781_551# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=0 ps=0
M1096 a_711_164# b2 a_699_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1097 gnd clk a_n124_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1098 a_853_889# cin vdd w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 a_817_551# a0 a_853_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 a_n131_15# clk vdd w_n139_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1101 a3 a_414_15# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1102 a_759_455# a0 vdd w_686_449# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1103 a_414_15# a_368_15# vdd w_406_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1104 gnd a0 a_690_n370# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1105 a_766_50# cin vdd w_693_44# CMOSP w=40 l=2
+  ad=600 pd=190 as=0 ps=0
M1106 a_709_551# a3 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1107 c3 a_711_164# vdd w_919_379# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1108 a_730_n123# b0 a_766_n123# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 a_n176_n239# b0_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1110 a_745_889# b2 a_733_889# w_692_883# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1111 gnd a2 a_745_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 a_n7_12# clk a_n7_96# w_n21_88# CMOSP w=80 l=2
+  ad=400 pd=170 as=800 ps=180
M1113 a_733_889# b2 a_781_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 a_699_455# a2 vdd w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 a_735_164# b1 a_723_164# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1116 b0 a_n86_n236# vdd w_n62_n160# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1117 b0 a_n86_n236# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1118 a_723_164# b1 a_771_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 gnd clk a_43_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 a1 a_83_15# vdd w_107_91# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1121 a_n124_15# a_n175_12# a_n131_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1122 a_730_50# b0 a_766_50# w_815_44# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 a_421_15# clk a_414_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1124 a_730_50# a0 a_766_50# w_693_44# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 a_718_50# a1 a_730_n123# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1126 a_158_n155# b2_in vdd w_144_n163# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1127 c1 n010 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1128 vdd a0 a_690_n308# w_677_n314# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 a_89_n236# clk a_82_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1130 a_n79_n236# clk a_n86_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1131 gnd a_368_15# a_421_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 cout a_721_551# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1133 a_829_551# b0 a_817_551# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1134 a_714_n370# cin gnd Gnd CMOSN w=20 l=2
+  ad=300 pd=110 as=0 ps=0
M1135 a_817_889# b1 a_781_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 a_323_n155# b3_in vdd w_309_n163# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1137 a_781_551# a1 a_817_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 a_n176_n239# clk a_n176_n155# w_n190_n163# CMOSP w=80 l=2
+  ad=400 pd=170 as=800 ps=180
M1139 a_817_889# a0 a_853_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 a_771_455# b0 a_759_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 a_807_164# a0 a_771_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 a_709_889# a3 vdd w_692_883# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1143 a_721_551# b3 a_709_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 a_718_50# a1 a_730_50# w_693_44# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 vdd a2 a_745_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 a_769_551# a1 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1147 gnd a1 a_735_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 a_413_n236# a_367_n236# vdd w_405_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1149 a_817_551# b0 a_853_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 n010 b0 a_714_n370# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 gnd a_n132_n236# a_n79_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 a_771_164# a1 a_723_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 a_374_n236# a_323_n239# a_367_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1154 a_706_n123# a_704_n129# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 a_771_455# b0 a_807_455# w_844_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1156 a_158_n239# clk a_158_n155# w_144_n163# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1157 gnd clk a_n125_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 a_721_551# a3 a_733_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 a0 a_n85_15# vdd w_n61_91# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1160 a_714_n308# cin vdd w_677_n314# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1161 gnd a_36_n236# a_89_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 a_n8_n239# b1_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1163 a2 a_249_15# vdd w_273_91# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1164 n010 a0 a_714_n370# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 b2 a_248_n236# vdd w_272_n160# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1166 a_711_164# a2 a_723_455# w_883_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 b2 a_248_n236# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1168 a_36_n236# clk vdd w_28_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1169 a_323_n239# clk a_323_n155# w_309_n163# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1170 a_n176_n155# b0_in vdd w_n190_n163# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 gnd a0 a_829_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 a_829_889# b0 a_817_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 b3 a_413_n236# vdd w_437_n160# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1174 c1 n010 vdd w_782_n313# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1175 b3 a_413_n236# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1176 a_781_889# a1 a_817_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 gnd cin a_807_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 a_721_551# b3 a_709_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 n010 b0 a_714_n308# w_749_n314# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1180 a_781_551# b1 a_769_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 a_n7_96# a1_in vdd w_n21_88# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 a_769_889# a1 vdd w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 a_711_164# b2 a_699_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a3 cin 0.32fF
C1 a_718_50# a0 0.13fF
C2 w_902_883# a_853_889# 0.06fF
C3 a1 b0 3.21fF
C4 b1 b0 7.24fF
C5 w_144_n163# vdd 0.20fF
C6 w_n61_91# vdd 0.06fF
C7 w_815_44# a_766_50# 0.06fF
C8 a_745_889# vdd 0.41fF
C9 w_692_883# a_829_889# 0.02fF
C10 a_n176_n239# b0_in 0.07fF
C11 b2 a_733_551# 0.21fF
C12 a_781_889# b0 0.10fF
C13 a0 a_716_n126# 0.15fF
C14 w_107_91# vdd 0.06fF
C15 a_374_n236# gnd 0.41fF
C16 a2 a1 5.36fF
C17 w_870_16# c2 0.06fF
C18 a2 b1 1.93fF
C19 b2 w_686_449# 0.13fF
C20 a_n79_n236# gnd 0.41fF
C21 a_36_n236# a_43_n236# 0.41fF
C22 a_730_n123# a0 0.13fF
C23 w_902_883# b0 0.06fF
C24 a_721_551# cin 0.17fF
C25 a_733_889# a0 0.15fF
C26 w_75_90# vdd 0.17fF
C27 a_413_n236# a_367_n236# 0.54fF
C28 gnd c2 0.21fF
C29 a3 gnd 0.21fF
C30 a_781_889# a2 0.10fF
C31 b0_in w_n190_n163# 0.08fF
C32 w_686_449# a_735_455# 0.02fF
C33 w_359_n161# vdd 0.17fF
C34 a_202_n236# w_194_n161# 0.10fF
C35 a_853_889# a0 0.09fF
C36 w_692_883# a1 0.13fF
C37 a_706_50# vdd 0.41fF
C38 w_692_883# b1 0.13fF
C39 a_704_n129# cin 0.08fF
C40 w_692_883# a_709_889# 0.02fF
C41 a_n176_n239# gnd 0.44fF
C42 a_781_551# cin 0.09fF
C43 a_718_50# w_693_44# 0.09fF
C44 a_771_455# b0 0.01fF
C45 a_n86_n236# b0 0.05fF
C46 b1_in a_n8_n239# 0.07fF
C47 a_n8_n239# vdd 0.03fF
C48 c1 n010 0.05fF
C49 a_781_889# w_692_883# 0.19fF
C50 a_n85_15# w_n93_90# 0.10fF
C51 a_413_n236# b3 0.05fF
C52 b2 a1 1.12fF
C53 a_n175_12# gnd 0.44fF
C54 b3 b0 0.69fF
C55 clk vdd 1.34fF
C56 b2 b1 6.06fF
C57 a_323_n155# vdd 0.89fF
C58 a_n131_15# clk 0.86fF
C59 a_n176_n155# vdd 0.88fF
C60 w_144_n163# a_158_n239# 0.11fF
C61 gnd a_721_551# 0.04fF
C62 a3 w_438_91# 0.06fF
C63 a_414_15# w_406_90# 0.10fF
C64 b0 a0 6.91fF
C65 a_367_n236# a_323_n239# 0.13fF
C66 a_817_889# a_829_889# 0.41fF
C67 a_n175_12# a_n175_96# 0.82fF
C68 n010 a_690_n308# 0.41fF
C69 a_n132_n236# clk 0.85fF
C70 b2 a_781_889# 0.10fF
C71 b0 a_723_455# 0.15fF
C72 a_n7_12# a_37_15# 0.13fF
C73 a_249_15# vdd 0.86fF
C74 c1 vdd 0.77fF
C75 w_686_449# vdd 0.17fF
C76 b3 a2 0.53fF
C77 a_829_889# vdd 0.41fF
C78 a2 a0 1.11fF
C79 a_36_n236# vdd 0.86fF
C80 vdd a_690_n308# 0.41fF
C81 a_90_15# gnd 0.41fF
C82 b3 w_692_883# 0.14fF
C83 a_817_889# a1 0.09fF
C84 a_368_15# a_324_12# 0.13fF
C85 a_414_15# vdd 0.86fF
C86 w_692_883# a0 0.13fF
C87 w_n94_n161# vdd 0.17fF
C88 vdd a_203_15# 0.86fF
C89 a_733_551# cin 0.10fF
C90 a1 vdd 0.89fF
C91 a_781_889# a_817_889# 1.20fF
C92 b1 vdd 0.81fF
C93 vdd a_709_889# 0.41fF
C94 b3 b2 4.09fF
C95 a_324_96# w_310_88# 0.02fF
C96 a_n132_n236# w_n94_n161# 0.07fF
C97 clk a_158_n239# 0.52fF
C98 a_807_455# vdd 0.41fF
C99 a_759_455# w_686_449# 0.02fF
C100 w_686_449# cin 0.06fF
C101 b2 a_248_n236# 0.05fF
C102 b0 w_693_44# 0.08fF
C103 gnd a_151_67# 0.02fF
C104 w_107_91# a_83_15# 0.08fF
C105 a_771_164# a1 0.01fF
C106 a_723_164# b0 0.15fF
C107 a_817_889# w_902_883# 0.06fF
C108 a_90_15# a_83_15# 0.41fF
C109 b2 a0 0.90fF
C110 w_n189_88# a0_in 0.08fF
C111 a_n86_n236# w_n62_n160# 0.08fF
C112 a_771_164# b1 0.01fF
C113 gnd a_n8_n239# 0.44fF
C114 w_749_n314# b0 0.10fF
C115 w_677_n314# a_690_n308# 0.02fF
C116 a_209_n236# a_202_n236# 0.41fF
C117 w_74_n161# a_82_n236# 0.10fF
C118 a_730_n123# a_766_n123# 0.41fF
C119 a_742_n123# a_754_n123# 0.21fF
C120 w_75_90# a_83_15# 0.10fF
C121 a_714_n308# a0 0.08fF
C122 a_723_455# a_735_455# 0.41fF
C123 a_n7_12# vdd 0.03fF
C124 gnd a_769_551# 0.21fF
C125 a_367_n236# vdd 0.86fF
C126 w_883_449# a2 0.06fF
C127 a1 cin 1.01fF
C128 a_420_n236# a_413_n236# 0.41fF
C129 a_249_15# gnd 0.10fF
C130 c1 gnd 0.23fF
C131 gnd a_853_551# 0.21fF
C132 a3 a_721_551# 0.24fF
C133 a0 n010 0.01fF
C134 b1 cin 0.67fF
C135 a_n86_n236# vdd 0.85fF
C136 cin a_807_455# 0.06fF
C137 a_255_n236# gnd 0.41fF
C138 w_n22_n163# a_n8_n239# 0.11fF
C139 a_817_889# a0 0.18fF
C140 a_781_889# cin 0.10fF
C141 w_n140_n161# clk 0.07fF
C142 a_n86_n236# a_n132_n236# 0.54fF
C143 clk a_83_15# 0.13fF
C144 a_202_n236# vdd 0.86fF
C145 a_n176_n239# w_n190_n163# 0.11fF
C146 b3 vdd 0.80fF
C147 gnd a_421_15# 0.41fF
C148 w_n22_n163# clk 0.08fF
C149 a_n7_96# a_n7_12# 0.82fF
C150 a_248_n236# vdd 0.86fF
C151 cout w_985_824# 0.06fF
C152 a0 vdd 2.07fF
C153 w_n189_88# vdd 0.20fF
C154 a_711_164# w_686_449# 0.03fF
C155 gnd a_414_15# 0.10fF
C156 w_815_44# b0 0.08fF
C157 a1 a_718_n123# 0.07fF
C158 w_272_n160# b2 0.06fF
C159 gnd a1 0.40fF
C160 w_360_90# vdd 0.17fF
C161 b1 a_718_n123# 0.03fF
C162 gnd b1 0.60fF
C163 a_771_164# a0 0.01fF
C164 a1_in gnd 0.02fF
C165 a_771_455# cin 0.01fF
C166 a_714_n308# w_749_n314# 0.06fF
C167 a_759_455# a_771_455# 0.41fF
C168 a_730_50# a1 0.06fF
C169 w_240_n161# a_202_n236# 0.07fF
C170 a_829_551# a_817_551# 0.21fF
C171 a_742_50# vdd 0.41fF
C172 b3 cin 2.05fF
C173 w_240_n161# a_248_n236# 0.10fF
C174 a_413_n236# w_437_n160# 0.08fF
C175 w_677_n314# a0 0.21fF
C176 a_711_164# a1 0.28fF
C177 w_749_n314# n010 0.06fF
C178 cout vdd 0.41fF
C179 a1 a_83_15# 0.05fF
C180 a_159_12# w_145_88# 0.11fF
C181 a_414_15# w_438_91# 0.08fF
C182 a_730_n123# a_718_50# 0.47fF
C183 a_256_15# gnd 0.41fF
C184 a_711_164# b1 0.36fF
C185 gnd a_89_n236# 0.41fF
C186 a0 cin 5.43fF
C187 a_324_12# a3_in 0.07fF
C188 a_n7_12# gnd 0.44fF
C189 a_n131_15# a_n124_15# 0.41fF
C190 cin a_723_455# 0.08fF
C191 a_817_551# b0 0.23fF
C192 a_202_n236# a_158_n239# 0.13fF
C193 w_693_44# vdd 0.10fF
C194 w_195_90# clk 0.07fF
C195 a_n86_n236# gnd 0.10fF
C196 a3 a_733_551# 1.49fF
C197 a_n176_n239# clk 0.52fF
C198 w_272_n160# vdd 0.06fF
C199 w_844_449# a_807_455# 0.06fF
C200 a_723_164# a_735_164# 0.21fF
C201 a_n176_n155# a_n176_n239# 0.82fF
C202 w_n139_90# clk 0.07fF
C203 a_771_164# a_723_164# 0.50fF
C204 gnd b3 0.30fF
C205 a_759_164# a_771_164# 0.21fF
C206 a_n175_12# clk 0.52fF
C207 gnd a_248_n236# 0.10fF
C208 a0 a_718_n123# 0.15fF
C209 clk w_310_88# 0.08fF
C210 gnd a0 0.61fF
C211 a_718_50# b0 0.20fF
C212 w_n190_n163# clk 0.08fF
C213 a_n176_n155# w_n190_n163# 0.02fF
C214 a_769_889# w_692_883# 0.02fF
C215 a_766_50# vdd 0.87fF
C216 a_721_551# a_733_551# 1.23fF
C217 cin w_693_44# 0.08fF
C218 a_367_n236# w_405_n161# 0.07fF
C219 a3 a_414_15# 0.05fF
C220 a_730_50# a0 0.13fF
C221 w_n189_88# a_n175_96# 0.02fF
C222 a_158_n155# vdd 0.89fF
C223 a_723_164# cin 0.08fF
C224 gnd a_n78_15# 0.41fF
C225 a3 a1 0.92fF
C226 b0 a_716_n126# 0.15fF
C227 a3 b1 0.64fF
C228 w_195_90# a_203_15# 0.10fF
C229 a_368_15# w_406_90# 0.07fF
C230 w_144_n163# clk 0.08fF
C231 a_771_455# w_844_449# 0.06fF
C232 w_782_n313# n010 0.08fF
C233 a_711_164# a0 0.26fF
C234 a_781_551# a_769_551# 0.21fF
C235 w_106_n160# b1 0.06fF
C236 a_733_551# a_781_551# 0.77fF
C237 a_711_164# a_723_455# 1.40fF
C238 w_241_90# vdd 0.17fF
C239 a_730_n123# b0 0.67fF
C240 a_853_551# a_781_551# 0.14fF
C241 a_733_889# b0 0.15fF
C242 cout gnd 0.21fF
C243 a_374_n236# a_367_n236# 0.41fF
C244 a_44_15# a_37_15# 0.41fF
C245 w_n93_90# vdd 0.17fF
C246 gnd a_n124_15# 0.41fF
C247 a_n131_15# w_n93_90# 0.07fF
C248 a_730_50# a_742_50# 0.41fF
C249 w_782_n313# vdd 0.10fF
C250 a_n85_15# vdd 0.85fF
C251 a_n131_15# a_n85_15# 0.54fF
C252 w_74_n161# vdd 0.17fF
C253 w_359_n161# clk 0.07fF
C254 a_721_551# a1 0.35fF
C255 a_733_889# a2 0.15fF
C256 w_309_n163# a_323_n239# 0.11fF
C257 w_28_n161# vdd 0.17fF
C258 a_759_164# gnd 0.21fF
C259 a_721_551# b1 0.25fF
C260 a_n86_n236# a_n79_n236# 0.41fF
C261 a_368_15# vdd 0.86fF
C262 a_721_551# a_709_889# 0.41fF
C263 a_733_889# w_941_883# 0.06fF
C264 a_375_15# a_368_15# 0.41fF
C265 a_n132_n236# a_n125_n236# 0.41fF
C266 a_730_50# w_693_44# 0.06fF
C267 clk a_n8_n239# 0.52fF
C268 a_704_n129# a1 0.09fF
C269 a2 w_273_91# 0.06fF
C270 w_437_n160# vdd 0.06fF
C271 a_781_551# a1 0.09fF
C272 a_699_455# vdd 0.41fF
C273 a_704_n129# b1 0.02fF
C274 a_733_889# w_692_883# 0.07fF
C275 a_781_551# b1 0.09fF
C276 a_158_n155# a_158_n239# 0.82fF
C277 a_324_12# vdd 0.03fF
C278 a_711_164# a_723_164# 0.96fF
C279 w_n21_88# vdd 0.20fF
C280 a3 b3 1.18fF
C281 w_107_91# a1 0.06fF
C282 a_769_889# vdd 0.41fF
C283 w_692_883# a_853_889# 0.03fF
C284 a_711_164# w_883_449# 0.06fF
C285 w_145_88# vdd 0.20fF
C286 a3 a0 0.93fF
C287 a_420_n236# gnd 0.41fF
C288 a_249_15# clk 0.13fF
C289 b2 a_733_889# 0.15fF
C290 a_36_n236# a_n8_n239# 0.13fF
C291 a2 b0 1.99fF
C292 gnd a_210_15# 0.41fF
C293 a_36_n236# clk 0.85fF
C294 a_766_50# a_730_50# 0.82fF
C295 a_766_n123# gnd 0.45fF
C296 a_n7_96# w_n21_88# 0.02fF
C297 b3 a_721_551# 0.17fF
C298 w_692_883# b0 0.06fF
C299 a_n175_12# w_n189_88# 0.11fF
C300 a_706_n123# a_718_n123# 0.21fF
C301 a_817_551# cin 0.12fF
C302 gnd a_706_n123# 0.21fF
C303 a_414_15# clk 0.13fF
C304 a_82_n236# vdd 0.86fF
C305 a_721_551# a0 0.25fF
C306 a_690_n370# n010 0.25fF
C307 clk a_203_15# 0.85fF
C308 a_n85_15# gnd 0.10fF
C309 w_815_44# a_730_50# 0.06fF
C310 w_309_n163# vdd 0.20fF
C311 w_692_883# a2 0.13fF
C312 gnd a_n125_n236# 0.41fF
C313 b2 b0 0.88fF
C314 a_733_551# a1 0.21fF
C315 a_704_n129# a0 0.15fF
C316 a_37_15# w_29_90# 0.10fF
C317 w_359_n161# a_367_n236# 0.10fF
C318 a_249_15# a_203_15# 0.54fF
C319 a_733_551# b1 0.21fF
C320 a_781_551# a0 0.18fF
C321 a_817_889# a_853_889# 1.79fF
C322 a_853_551# a1 0.09fF
C323 a1 w_686_449# 0.13fF
C324 w_n61_91# a0 0.06fF
C325 w_686_449# b1 0.13fF
C326 a_714_n370# n010 0.64fF
C327 b2 a2 3.61fF
C328 a_159_96# w_145_88# 0.02fF
C329 w_686_449# a_807_455# 0.03fF
C330 a_414_15# a_421_15# 0.41fF
C331 a_718_50# cin 0.06fF
C332 a_853_889# vdd 0.41fF
C333 w_n62_n160# b0 0.06fF
C334 gnd a_324_12# 0.44fF
C335 w_309_n163# b3_in 0.08fF
C336 cout a_721_551# 0.05fF
C337 a_n7_12# clk 0.52fF
C338 a_367_n236# clk 0.85fF
C339 w_273_91# vdd 0.06fF
C340 b0 n010 0.01fF
C341 w_194_n161# vdd 0.17fF
C342 a_159_12# vdd 0.03fF
C343 b2 w_692_883# 0.13fF
C344 a_249_15# a_256_15# 0.41fF
C345 a_n86_n236# clk 0.13fF
C346 a_817_889# b0 0.18fF
C347 cin a_716_n126# 0.08fF
C348 a_699_455# a_711_164# 0.41fF
C349 a1 b1 5.31fF
C350 a_413_n236# vdd 0.86fF
C351 a_718_50# w_870_16# 0.08fF
C352 a_202_n236# clk 0.85fF
C353 a_730_n123# cin 0.06fF
C354 b0 vdd 0.82fF
C355 a_733_889# cin 0.08fF
C356 a_718_50# a_718_n123# 0.01fF
C357 c3 vdd 0.41fF
C358 clk a_248_n236# 0.13fF
C359 a_771_455# w_686_449# 0.06fF
C360 a_718_50# gnd 0.04fF
C361 a_44_15# gnd 0.41fF
C362 a_781_889# a1 0.10fF
C363 a_781_889# b1 0.10fF
C364 w_n189_88# clk 0.08fF
C365 a_754_n123# a_766_n123# 0.21fF
C366 a_771_164# b0 0.01fF
C367 gnd a_82_n236# 0.10fF
C368 a_733_551# a0 0.21fF
C369 a2 vdd 0.84fF
C370 a_718_50# a_730_50# 1.84fF
C371 clk w_360_90# 0.07fF
C372 w_29_90# vdd 0.17fF
C373 a_853_551# a0 0.09fF
C374 a_255_n236# a_248_n236# 0.41fF
C375 a_817_889# w_692_883# 0.11fF
C376 w_686_449# a0 0.13fF
C377 w_686_449# a_723_455# 0.06fF
C378 a_324_96# a_324_12# 0.82fF
C379 b2_in a_158_n239# 0.07fF
C380 a1_in a_n7_12# 0.07fF
C381 a_730_n123# a_718_n123# 0.21fF
C382 a_323_n239# vdd 0.03fF
C383 a_n86_n236# w_n94_n161# 0.10fF
C384 w_677_n314# b0 0.10fF
C385 a_771_455# a1 0.01fF
C386 w_692_883# vdd 0.14fF
C387 a_37_15# vdd 0.86fF
C388 a_690_n370# gnd 0.21fF
C389 a_706_50# w_693_44# 0.02fF
C390 a_771_455# b1 0.01fF
C391 b0 cin 1.69fF
C392 a_n8_n155# vdd 0.89fF
C393 a_159_12# a_159_96# 0.82fF
C394 a_771_455# a_807_455# 1.04fF
C395 a_714_n308# n010 1.06fF
C396 b3 a1 0.77fF
C397 gnd b2_in 0.02fF
C398 gnd a_745_551# 0.21fF
C399 a_158_n155# w_144_n163# 0.02fF
C400 b3 b1 0.60fF
C401 b2 vdd 0.84fF
C402 a2 cin 0.59fF
C403 a1 a0 8.37fF
C404 a_159_12# gnd 0.44fF
C405 gnd a_829_551# 0.21fF
C406 a1 a_723_455# 0.15fF
C407 b3_in a_323_n239# 0.07fF
C408 b1 a0 1.31fF
C409 gnd a_714_n370# 0.21fF
C410 b1 a_723_455# 0.15fF
C411 a_735_455# vdd 0.41fF
C412 w_919_379# c3 0.06fF
C413 a_714_n308# vdd 0.41fF
C414 w_985_824# vdd 0.06fF
C415 gnd a3_in 0.02fF
C416 a_781_889# a0 0.21fF
C417 a_413_n236# gnd 0.10fF
C418 w_406_90# vdd 0.17fF
C419 b0 a_718_n123# 0.18fF
C420 gnd b0 1.09fF
C421 w_692_883# cin 0.06fF
C422 w_n62_n160# vdd 0.06fF
C423 gnd c3 0.21fF
C424 a_n85_15# w_n61_91# 0.08fF
C425 vdd n010 0.39fF
C426 a_324_12# w_310_88# 0.11fF
C427 a_718_50# c2 0.05fF
C428 a_730_50# b0 0.13fF
C429 gnd a2 0.41fF
C430 b2 cin 0.47fF
C431 a_711_164# b0 0.26fF
C432 a_714_n308# w_677_n314# 0.03fF
C433 a_771_455# a0 0.01fF
C434 w_106_n160# a_82_n236# 0.08fF
C435 a_711_164# c3 0.05fF
C436 a_781_551# a_817_551# 0.83fF
C437 a_771_455# a_723_455# 0.97fF
C438 a1 w_693_44# 0.15fF
C439 a_202_n236# a_248_n236# 0.54fF
C440 a_n131_15# vdd 0.85fF
C441 gnd a_323_n239# 0.44fF
C442 a_723_164# a1 0.15fF
C443 b1 w_693_44# 0.15fF
C444 a_723_164# b1 0.15fF
C445 b3 a0 0.69fF
C446 a_n132_n236# vdd 0.85fF
C447 a_413_n236# w_405_n161# 0.10fF
C448 a_711_164# a2 0.26fF
C449 w_677_n314# n010 0.34fF
C450 w_844_449# b0 0.06fF
C451 gnd a_43_n236# 0.41fF
C452 cin n010 0.00fF
C453 a0 a_723_455# 0.15fF
C454 gnd a0_in 0.02fF
C455 a_249_15# w_241_90# 0.10fF
C456 gnd b2 0.62fF
C457 a_730_n123# a_742_n123# 0.21fF
C458 a_n85_15# clk 0.13fF
C459 a_n7_96# vdd 0.89fF
C460 a_817_889# cin 0.09fF
C461 gnd a_709_551# 0.21fF
C462 a_37_15# a_83_15# 0.54fF
C463 w_28_n161# clk 0.07fF
C464 w_677_n314# vdd 0.03fF
C465 a_368_15# clk 0.85fF
C466 w_240_n161# vdd 0.17fF
C467 w_782_n313# c1 0.06fF
C468 a_759_455# vdd 0.41fF
C469 cin vdd 0.34fF
C470 a_210_15# a_203_15# 0.41fF
C471 a_n8_n155# w_n22_n163# 0.02fF
C472 a_209_n236# gnd 0.41fF
C473 w_145_88# a_151_67# 0.08fF
C474 a_721_551# a_733_889# 1.48fF
C475 a_711_164# b2 0.18fF
C476 a_771_164# cin 0.01fF
C477 gnd n010 0.26fF
C478 w_74_n161# a_36_n236# 0.07fF
C479 a_158_n239# vdd 0.03fF
C480 a3 b0 1.72fF
C481 w_241_90# a_203_15# 0.07fF
C482 w_n21_88# clk 0.08fF
C483 clk a_324_12# 0.52fF
C484 w_28_n161# a_36_n236# 0.10fF
C485 a_159_96# vdd 0.89fF
C486 w_919_379# vdd 0.06fF
C487 a_699_455# w_686_449# 0.02fF
C488 w_145_88# clk 0.08fF
C489 a0 w_693_44# 0.15fF
C490 a_853_551# a_817_551# 0.78fF
C491 w_870_16# vdd 0.06fF
C492 a_706_50# a_718_50# 0.41fF
C493 a_723_164# a0 0.15fF
C494 w_272_n160# a_248_n236# 0.08fF
C495 a_745_889# a_733_889# 0.41fF
C496 a3 a2 2.78fF
C497 w_677_n314# cin 0.10fF
C498 b1_in gnd 0.02fF
C499 w_310_88# a3_in 0.08fF
C500 a_414_15# a_368_15# 0.54fF
C501 a3 w_941_883# 0.06fF
C502 a_375_15# gnd 0.41fF
C503 w_883_449# a_723_455# 0.06fF
C504 w_144_n163# b2_in 0.08fF
C505 a_771_164# a_807_164# 0.50fF
C506 gnd a_735_164# 0.21fF
C507 a_721_551# b0 0.25fF
C508 a_n175_96# vdd 0.88fF
C509 a3 w_692_883# 0.06fF
C510 a_742_50# w_693_44# 0.02fF
C511 clk a_82_n236# 0.13fF
C512 a_817_551# a1 0.12fF
C513 a_704_n129# b0 0.08fF
C514 w_n140_n161# vdd 0.17fF
C515 a_83_15# vdd 0.86fF
C516 gnd b3_in 0.02fF
C517 a_781_551# b0 0.09fF
C518 w_309_n163# clk 0.08fF
C519 b1_in w_n22_n163# 0.08fF
C520 w_309_n163# a_323_n155# 0.02fF
C521 a_721_551# a2 0.32fF
C522 w_n22_n163# vdd 0.20fF
C523 a_807_164# cin 0.09fF
C524 a3 b2 0.65fF
C525 a_n132_n236# w_n140_n161# 0.10fF
C526 w_438_91# vdd 0.06fF
C527 a_721_551# w_941_883# 0.06fF
C528 a1_in w_n21_88# 0.08fF
C529 cin a_718_n123# 0.07fF
C530 gnd b0_in 0.02fF
C531 a_781_889# a_769_889# 0.41fF
C532 w_405_n161# vdd 0.17fF
C533 a_781_551# a2 0.09fF
C534 a_36_n236# a_82_n236# 0.54fF
C535 a_721_551# w_692_883# 0.03fF
C536 a_159_12# a_151_67# 0.07fF
C537 gnd a_699_164# 0.21fF
C538 a_730_50# cin 0.06fF
C539 a_324_96# vdd 0.89fF
C540 gnd a_158_n239# 0.44fF
C541 a_n175_12# a0_in 0.07fF
C542 a_718_50# a1 0.06fF
C543 a_n7_12# w_n21_88# 0.11fF
C544 w_194_n161# clk 0.07fF
C545 a_718_50# b1 0.09fF
C546 a_733_551# a_745_551# 0.21fF
C547 a_711_164# cin 0.19fF
C548 a_159_12# clk 0.52fF
C549 a_n85_15# a0 0.05fF
C550 b2 a_721_551# 0.41fF
C551 gnd a_807_164# 0.23fF
C552 a_745_889# w_692_883# 0.02fF
C553 a_249_15# w_273_91# 0.08fF
C554 a_721_551# a_709_551# 0.21fF
C555 a_82_n236# b1 0.05fF
C556 a_711_164# a_699_164# 0.21fF
C557 a_766_50# w_693_44# 0.03fF
C558 b3 w_437_n160# 0.06fF
C559 a_413_n236# clk 0.13fF
C560 a1 a_716_n126# 0.08fF
C561 a_721_551# w_985_824# 0.08fF
C562 b1 a_716_n126# 0.04fF
C563 b2 a_781_551# 0.09fF
C564 a_368_15# w_360_90# 0.10fF
C565 vdd c2 0.41fF
C566 a_n85_15# a_n78_15# 0.41fF
C567 a3 vdd 0.80fF
C568 a_711_164# w_919_379# 0.08fF
C569 w_106_n160# vdd 0.06fF
C570 a_37_15# w_75_90# 0.07fF
C571 a_733_551# b0 0.21fF
C572 a_817_551# a0 0.23fF
C573 a_730_n123# a1 0.06fF
C574 a_733_889# a1 0.15fF
C575 w_195_90# vdd 0.17fF
C576 a_733_889# b1 0.15fF
C577 a_n176_n239# vdd 0.03fF
C578 a_82_n236# a_89_n236# 0.41fF
C579 w_686_449# b0 0.06fF
C580 a_853_889# a1 0.09fF
C581 a_711_164# gnd 0.04fF
C582 w_n139_90# vdd 0.17fF
C583 gnd a_83_15# 0.10fF
C584 a_n131_15# w_n139_90# 0.10fF
C585 clk w_29_90# 0.07fF
C586 a_781_889# a_733_889# 1.27fF
C587 a_n132_n236# a_n176_n239# 0.13fF
C588 a_733_551# a2 0.21fF
C589 a_n175_12# vdd 0.03fF
C590 a_n131_15# a_n175_12# 0.13fF
C591 a_159_12# a_203_15# 0.13fF
C592 w_310_88# vdd 0.20fF
C593 a_n8_n155# a_n8_n239# 0.82fF
C594 a_249_15# a2 0.05fF
C595 a_781_889# a_853_889# 0.16fF
C596 clk a_323_n239# 0.52fF
C597 a2 w_686_449# 0.06fF
C598 a_323_n155# a_323_n239# 0.82fF
C599 w_n190_n163# vdd 0.20fF
C600 a_37_15# clk 0.85fF
C601 a_714_n370# Gnd 0.13fF
C602 a_690_n370# Gnd 0.04fF
C603 c1 Gnd 0.14fF
C604 a_714_n308# Gnd 0.15fF
C605 a_690_n308# Gnd 0.00fF
C606 n010 Gnd 3.19fF
C607 a_420_n236# Gnd 0.02fF
C608 a_374_n236# Gnd 0.02fF
C609 a_255_n236# Gnd 0.02fF
C610 a_209_n236# Gnd 0.02fF
C611 a_766_n123# Gnd 0.29fF
C612 a_754_n123# Gnd 0.02fF
C613 a_742_n123# Gnd 0.02fF
C614 a_730_n123# Gnd 0.49fF
C615 a_718_n123# Gnd 0.53fF
C616 a_706_n123# Gnd 0.02fF
C617 c2 Gnd 0.11fF
C618 a_716_n126# Gnd 0.53fF
C619 a_704_n129# Gnd 0.55fF
C620 a_413_n236# Gnd 0.75fF
C621 a_323_n239# Gnd 0.48fF
C622 a_323_n155# Gnd 0.00fF
C623 a_89_n236# Gnd 0.02fF
C624 a_43_n236# Gnd 0.02fF
C625 a_248_n236# Gnd 0.75fF
C626 a_158_n239# Gnd 0.48fF
C627 a_158_n155# Gnd 0.00fF
C628 a_n79_n236# Gnd 0.02fF
C629 a_n125_n236# Gnd 0.02fF
C630 a_82_n236# Gnd 0.75fF
C631 a_n8_n239# Gnd 0.48fF
C632 a_n8_n155# Gnd 0.00fF
C633 a_n86_n236# Gnd 0.75fF
C634 a_n176_n239# Gnd 0.48fF
C635 a_n176_n155# Gnd 0.00fF
C636 a_367_n236# Gnd 1.01fF
C637 b3_in Gnd 0.21fF
C638 a_202_n236# Gnd 1.01fF
C639 b2_in Gnd 0.34fF
C640 a_36_n236# Gnd 1.01fF
C641 b1_in Gnd 0.15fF
C642 a_n132_n236# Gnd 1.01fF
C643 b0_in Gnd 0.15fF
C644 a_766_50# Gnd 0.18fF
C645 a_742_50# Gnd 0.00fF
C646 a_730_50# Gnd 0.47fF
C647 a_718_50# Gnd 2.46fF
C648 a_706_50# Gnd 0.00fF
C649 a_421_15# Gnd 0.02fF
C650 a_375_15# Gnd 0.02fF
C651 a_256_15# Gnd 0.02fF
C652 a_210_15# Gnd 0.02fF
C653 a_807_164# Gnd 0.22fF
C654 a_771_164# Gnd 1.17fF
C655 a_759_164# Gnd 0.02fF
C656 a_735_164# Gnd 0.02fF
C657 a_723_164# Gnd 1.01fF
C658 a_699_164# Gnd 0.02fF
C659 a_414_15# Gnd 0.75fF
C660 a_324_12# Gnd 0.25fF
C661 a_324_96# Gnd 0.00fF
C662 a_90_15# Gnd 0.02fF
C663 a_44_15# Gnd 0.02fF
C664 a_249_15# Gnd 0.75fF
C665 a_159_96# Gnd 0.00fF
C666 a_n78_15# Gnd 0.02fF
C667 a_n124_15# Gnd 0.02fF
C668 a_83_15# Gnd 0.75fF
C669 a_n7_12# Gnd 0.18fF
C670 a_n7_96# Gnd 0.00fF
C671 a_n85_15# Gnd 0.75fF
C672 a_n175_12# Gnd 0.18fF
C673 a_n175_96# Gnd 0.00fF
C674 a_368_15# Gnd 1.01fF
C675 a3_in Gnd 0.34fF
C676 a_203_15# Gnd 1.01fF
C677 a_151_67# Gnd 0.34fF
C678 a_37_15# Gnd 1.01fF
C679 a1_in Gnd 0.28fF
C680 a_n131_15# Gnd 1.01fF
C681 clk Gnd 0.09fF
C682 a0_in Gnd 0.28fF
C683 c3 Gnd 0.10fF
C684 a_807_455# Gnd 0.20fF
C685 a_771_455# Gnd 1.16fF
C686 a_759_455# Gnd 0.00fF
C687 a_735_455# Gnd 0.00fF
C688 a_723_455# Gnd 0.92fF
C689 a_711_164# Gnd 3.38fF
C690 a_699_455# Gnd 0.00fF
C691 a_853_551# Gnd 0.30fF
C692 a_829_551# Gnd 0.02fF
C693 a_817_551# Gnd 0.89fF
C694 a_781_551# Gnd 1.29fF
C695 a_769_551# Gnd 0.02fF
C696 a_745_551# Gnd 0.02fF
C697 a_733_551# Gnd 2.00fF
C698 a_709_551# Gnd 0.02fF
C699 gnd Gnd 19.56fF
C700 cout Gnd 0.10fF
C701 a_853_889# Gnd 0.23fF
C702 a_829_889# Gnd 0.00fF
C703 a_817_889# Gnd 0.59fF
C704 a_781_889# Gnd 0.98fF
C705 a_769_889# Gnd 0.00fF
C706 a_745_889# Gnd 0.00fF
C707 a_733_889# Gnd 1.46fF
C708 a_721_551# Gnd 4.42fF
C709 a_709_889# Gnd 0.00fF
C710 vdd Gnd 17.67fF
C711 cin Gnd 16.57fF
C712 a0 Gnd 33.77fF
C713 b0 Gnd 33.73fF
C714 b1 Gnd 28.22fF
C715 a1 Gnd 30.63fF
C716 a2 Gnd 26.32fF
C717 b2 Gnd 24.26fF
C718 b3 Gnd 16.47fF
C719 a3 Gnd 18.74fF
C720 w_782_n313# Gnd 1.25fF
C721 w_749_n314# Gnd 1.38fF
C722 w_677_n314# Gnd 3.51fF
C723 w_437_n160# Gnd 1.46fF
C724 w_405_n161# Gnd 2.53fF
C725 w_359_n161# Gnd 2.53fF
C726 w_309_n163# Gnd 3.68fF
C727 w_272_n160# Gnd 1.46fF
C728 w_240_n161# Gnd 2.53fF
C729 w_194_n161# Gnd 2.53fF
C730 w_144_n163# Gnd 0.01fF
C731 w_106_n160# Gnd 1.46fF
C732 w_74_n161# Gnd 2.53fF
C733 w_28_n161# Gnd 2.53fF
C734 w_n22_n163# Gnd 3.68fF
C735 w_n62_n160# Gnd 1.46fF
C736 w_n94_n161# Gnd 2.53fF
C737 w_n140_n161# Gnd 2.53fF
C738 w_n190_n163# Gnd 3.68fF
C739 w_870_16# Gnd 1.25fF
C740 w_815_44# Gnd 1.25fF
C741 w_693_44# Gnd 5.64fF
C742 w_438_91# Gnd 1.46fF
C743 w_406_90# Gnd 2.53fF
C744 w_360_90# Gnd 2.53fF
C745 w_310_88# Gnd 0.04fF
C746 w_273_91# Gnd 1.46fF
C747 w_241_90# Gnd 2.53fF
C748 w_195_90# Gnd 2.53fF
C749 w_145_88# Gnd 3.68fF
C750 w_107_91# Gnd 1.46fF
C751 w_75_90# Gnd 2.53fF
C752 w_29_90# Gnd 2.53fF
C753 w_n21_88# Gnd 3.68fF
C754 w_n61_91# Gnd 1.46fF
C755 w_n93_90# Gnd 2.53fF
C756 w_n139_90# Gnd 2.53fF
C757 w_n189_88# Gnd 3.68fF
C758 w_919_379# Gnd 1.25fF
C759 w_883_449# Gnd 1.33fF
C760 w_844_449# Gnd 1.33fF
C761 w_686_449# Gnd 7.72fF
C762 w_985_824# Gnd 1.25fF
C763 w_941_883# Gnd 1.33fF
C764 w_902_883# Gnd 1.33fF
C765 w_692_883# Gnd 10.49fF


.tran 10n 1u

.control
set hcopypscolor = 1 
set color0=white
set color1=black
run

*plot V(a0) V(b0)+2 V(cin)+4 V(c1)+6
*plot V(a1) V(b1)+2 V(c1)+4 V(c2)+6
plot V(a0) V(b0)+2 V(a1)+4 V(b1)+6
plot V(a2) V(b2)+2 V(c3)+4
*plot V(a0) V(b0)+2 V(a1)+4 V(b1)+6 
*plot V(a2) V(b2)+2 V(a3)+4 V(b3)+6 V(cout)+8
*plot V(a3) V(b3)+2 V(cout)+4
.endc
.end