magic
tech scmos
timestamp 1732053661
<< nwell >>
rect 115 82 228 135
rect 234 82 260 135
rect 132 81 169 82
rect 349 54 373 106
<< ntransistor >>
rect 137 24 139 44
rect 149 24 151 44
rect 161 24 163 44
rect 173 24 175 44
rect 185 24 187 44
rect 197 24 199 44
rect 209 24 211 44
rect 246 24 248 44
rect 360 23 362 43
<< ptransistor >>
rect 137 88 139 128
rect 149 88 151 128
rect 161 88 163 128
rect 173 88 175 128
rect 185 88 187 128
rect 197 88 199 128
rect 209 88 211 128
rect 246 88 248 128
rect 360 60 362 100
<< ndiffusion >>
rect 136 24 137 44
rect 139 24 140 44
rect 148 24 149 44
rect 151 24 152 44
rect 160 24 161 44
rect 163 24 164 44
rect 172 24 173 44
rect 175 24 176 44
rect 184 24 185 44
rect 187 24 188 44
rect 196 24 197 44
rect 199 24 200 44
rect 208 24 209 44
rect 211 24 212 44
rect 245 24 246 44
rect 248 24 249 44
rect 359 23 360 43
rect 362 23 363 43
<< pdiffusion >>
rect 136 88 137 128
rect 139 88 140 128
rect 148 88 149 128
rect 151 88 161 128
rect 163 88 173 128
rect 175 88 176 128
rect 184 88 185 128
rect 187 88 188 128
rect 196 88 197 128
rect 199 88 200 128
rect 208 88 209 128
rect 211 88 212 128
rect 245 88 246 128
rect 248 88 249 128
rect 359 60 360 100
rect 362 60 363 100
<< ndcontact >>
rect 132 24 136 44
rect 140 24 148 44
rect 152 24 160 44
rect 164 24 172 44
rect 176 24 184 44
rect 188 24 196 44
rect 200 24 208 44
rect 212 24 216 44
rect 241 24 245 44
rect 249 24 253 44
rect 355 23 359 43
rect 363 23 367 43
<< pdcontact >>
rect 132 88 136 128
rect 140 88 148 128
rect 176 88 184 128
rect 188 88 196 128
rect 200 88 208 128
rect 212 88 216 128
rect 241 88 245 128
rect 249 88 253 128
rect 355 60 359 100
rect 363 60 367 100
<< polysilicon >>
rect 137 128 139 131
rect 149 128 151 131
rect 161 128 163 131
rect 173 128 175 131
rect 185 128 187 131
rect 197 128 199 131
rect 209 128 211 131
rect 246 128 248 131
rect 360 100 362 106
rect 137 44 139 88
rect 149 44 151 88
rect 161 44 163 88
rect 173 44 175 88
rect 185 44 187 88
rect 197 44 199 88
rect 209 44 211 88
rect 246 44 248 88
rect 360 43 362 60
rect 137 19 139 24
rect 149 19 151 24
rect 161 20 163 24
rect 173 19 175 24
rect 185 19 187 24
rect 197 20 199 24
rect 209 20 211 24
rect 246 20 248 24
rect 360 19 362 23
<< polycontact >>
rect 136 131 140 135
rect 148 131 152 135
rect 160 131 164 135
rect 172 131 176 135
rect 184 131 188 135
rect 196 131 200 135
rect 208 131 212 135
rect 245 131 249 135
rect 355 47 360 51
<< metal1 >>
rect 152 88 160 128
rect 164 88 172 128
rect 216 93 221 97
rect 132 72 136 88
rect 154 72 158 88
rect 168 69 172 88
rect 190 72 194 88
rect 202 79 205 88
rect 242 79 245 88
rect 202 75 245 79
rect 349 106 373 110
rect 132 44 136 50
rect 168 44 172 64
rect 249 68 253 88
rect 355 100 359 106
rect 249 51 253 63
rect 363 51 367 60
rect 249 47 278 51
rect 339 47 355 51
rect 363 47 383 51
rect 249 44 253 47
rect 216 31 220 35
rect 132 16 136 24
rect 154 16 158 24
rect 168 4 172 24
rect 190 10 194 24
rect 202 14 206 24
rect 241 14 245 24
rect 202 10 245 14
rect 363 43 367 47
rect 249 5 253 24
rect 355 19 360 23
rect 349 15 373 19
<< m2contact >>
rect 221 93 227 98
rect 166 64 172 69
rect 249 63 255 68
rect 220 30 225 37
rect 168 -2 173 4
rect 248 -2 255 5
<< metal2 >>
rect 136 131 140 141
rect 148 131 152 143
rect 160 131 164 143
rect 172 131 176 141
rect 184 131 188 145
rect 196 131 200 153
rect 208 131 212 145
rect 245 131 249 141
rect 221 67 226 93
rect 172 64 249 67
rect 220 3 224 30
rect 173 -1 248 3
<< labels >>
rlabel metal1 192 13 192 13 1 gnd
rlabel metal2 247 137 247 137 5 b0
rlabel metal2 174 137 174 137 5 b0
rlabel metal2 186 137 186 137 5 a0
rlabel metal2 198 137 198 137 5 cin
rlabel metal2 210 137 210 137 5 a0
rlabel metal1 192 74 192 74 1 vdd
rlabel metal1 360 108 360 108 5 vdd
rlabel metal1 360 17 360 17 1 gnd
rlabel space 135 135 140 139 1 a1
rlabel space 148 135 153 139 1 b1
rlabel space 160 135 165 139 1 b1
rlabel metal1 132 72 136 79 1 vdd
<< end >>
