* SPICE3 file created from carry_one.ext - technology: scmos
.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY = 1.8
.param LAMBDA=0.09u
.global gnd vdd
Vdd vdd gnd 'SUPPLY'

V1 A0 gnd dc 0
V2 B0 gnd dc 'SUPPLY'
V3 cin gnd dc 'SUPPLY'
V4 A1 gnd dc 'SUPPLY'
V5 B1 gnd dc 'SUPPLY'

M1000 a_362_87# a1 vdd w_349_81# CMOSP w=120 l=2
+  ad=1200 pd=260 as=2000 ps=600
M1001 a_410_n117# a0 a_398_n117# Gnd CMOSN w=60 l=2
+  ad=600 pd=140 as=600 ps=140
M1002 a_362_n117# a_360_n125# gnd Gnd CMOSN w=60 l=2
+  ad=600 pd=140 as=400 ps=180
M1003 c2 a_374_87# vdd w_568_53# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1004 a_386_n117# a0 a_422_n117# Gnd CMOSN w=60 l=2
+  ad=1505 pd=412 as=905 ps=272
M1005 a_374_87# b1 a_362_87# w_349_81# CMOSP w=120 l=2
+  ad=1800 pd=510 as=0 ps=0
M1006 a_386_87# b1 a_374_87# w_349_81# CMOSP w=120 l=2
+  ad=3000 pd=770 as=0 ps=0
M1007 a_374_n117# a_372_n125# a_362_n117# Gnd CMOSN w=60 l=2
+  ad=600 pd=140 as=0 ps=0
M1008 a_374_87# a1 a_386_n117# Gnd CMOSN w=60 l=2
+  ad=300 pd=130 as=0 ps=0
M1009 a_398_87# b0 a_386_87# w_349_81# CMOSP w=120 l=2
+  ad=1200 pd=260 as=0 ps=0
M1010 a_386_n117# b1 a_374_n117# Gnd CMOSN w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 c2 a_374_87# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1012 a_398_n117# b0 a_386_n117# Gnd CMOSN w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 a_386_87# b0 a_422_87# w_471_81# CMOSP w=120 l=2
+  ad=0 pd=0 as=1800 ps=510
M1014 a_386_n117# b0 a_422_n117# Gnd CMOSN w=61 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 vdd a0 a_398_87# w_349_81# CMOSP w=120 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 a_422_87# cin vdd w_349_81# CMOSP w=120 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 a_386_87# a0 a_422_87# w_349_81# CMOSP w=120 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 a_374_87# a1 a_386_87# w_349_81# CMOSP w=120 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 a_422_n117# cin a_410_n117# Gnd CMOSN w=60 l=2
+  ad=0 pd=0 as=0 ps=0
C0 b0 a_386_87# 0.13fF
C1 a1 b0 1.18fF
C2 b1 a_374_87# 0.09fF
C3 b0 cin 0.24fF
C4 b0 a_386_n117# 0.67fF
C5 a0 a_374_n117# 0.15fF
C6 vdd a_362_87# 1.24fF
C7 a1 a_374_n117# 0.07fF
C8 b0 a_372_n125# 0.15fF
C9 a_374_87# c2 0.05fF
C10 cin a_374_n117# 0.07fF
C11 a_374_n117# a_386_n117# 0.62fF
C12 a_362_n117# a_374_n117# 0.62fF
C13 gnd a_362_n117# 0.62fF
C14 w_471_81# a_422_87# 0.15fF
C15 b0 w_471_81# 0.06fF
C16 a0 w_349_81# 0.13fF
C17 w_349_81# a_386_87# 0.06fF
C18 a_374_87# w_568_53# 0.08fF
C19 b1 a_360_n125# 0.02fF
C20 a1 w_349_81# 0.13fF
C21 a_386_87# a_398_87# 1.24fF
C22 b1 a0 0.15fF
C23 a_362_87# w_349_81# 0.02fF
C24 a_422_n117# a_386_n117# 1.25fF
C25 cin w_349_81# 0.06fF
C26 a0 a_374_87# 0.13fF
C27 a_374_87# a_386_87# 3.49fF
C28 vdd a_422_87# 1.70fF
C29 a1 b1 0.57fF
C30 c2 w_568_53# 0.06fF
C31 a1 a_374_87# 0.06fF
C32 b1 cin 0.08fF
C33 a_362_87# a_374_87# 1.24fF
C34 b0 a_374_n117# 0.18fF
C35 cin a_374_87# 0.06fF
C36 a_374_87# a_386_n117# 0.83fF
C37 b1 a_372_n125# 0.04fF
C38 a_386_n117# a_398_n117# 0.62fF
C39 w_349_81# a_422_87# 0.03fF
C40 a0 a_360_n125# 0.15fF
C41 b0 w_349_81# 0.06fF
C42 a1 a_360_n125# 0.09fF
C43 a0 a_386_87# 0.13fF
C44 a_422_n117# a_410_n117# 0.62fF
C45 b1 b0 0.48fF
C46 a1 a0 1.18fF
C47 vdd w_349_81# 0.18fF
C48 a1 a_386_87# 0.06fF
C49 cin a_360_n125# 0.08fF
C50 b0 a_374_87# 0.20fF
C51 vdd a_398_87# 1.24fF
C52 a_422_n117# gnd 0.45fF
C53 a0 cin 1.61fF
C54 cin a_386_87# 0.06fF
C55 a0 a_386_n117# 0.13fF
C56 a1 cin 0.17fF
C57 b1 a_374_n117# 0.03fF
C58 a1 a_386_n117# 0.06fF
C59 a0 a_372_n125# 0.15fF
C60 a_374_87# a_374_n117# 0.01fF
C61 a_398_n117# a_410_n117# 0.62fF
C62 a_374_87# gnd 0.04fF
C63 cin a_386_n117# 0.06fF
C64 a1 a_372_n125# 0.08fF
C65 vdd c2 0.41fF
C66 cin a_372_n125# 0.08fF
C67 c2 gnd 0.21fF
C68 w_471_81# a_386_87# 0.14fF
C69 w_349_81# a_398_87# 0.02fF
C70 b0 a_360_n125# 0.08fF
C71 b1 w_349_81# 0.13fF
C72 a_386_87# a_422_87# 2.47fF
C73 b0 a0 1.22fF
C74 a_374_87# w_349_81# 0.17fF
C75 vdd w_568_53# 0.06fF
C76 a_422_n117# Gnd 0.29fF
C77 a_410_n117# Gnd 0.02fF
C78 a_398_n117# Gnd 0.02fF
C79 a_386_n117# Gnd 0.49fF
C80 a_374_n117# Gnd 0.50fF
C81 a_362_n117# Gnd 0.02fF
C82 gnd Gnd 1.46fF
C83 c2 Gnd 0.11fF
C84 a_372_n125# Gnd 0.50fF
C85 a_360_n125# Gnd 0.50fF
C86 a_422_87# Gnd 0.17fF
C87 a_398_87# Gnd 0.00fF
C88 a_386_87# Gnd 0.47fF
C89 a_374_87# Gnd 2.63fF
C90 a_362_87# Gnd 0.00fF
C91 vdd Gnd 1.13fF
C92 cin Gnd 1.16fF
C93 a0 Gnd 2.47fF
C94 b0 Gnd 2.67fF
C95 b1 Gnd 1.50fF
C96 a1 Gnd 2.23fF
C97 w_568_53# Gnd 1.25fF
C98 w_471_81# Gnd 3.34fF
C99 w_349_81# Gnd 14.56fF

.tran 0.1n 1u

.control
set hcopypscolor = 1 
set color0=white
set color1=black
run

plot V(a0) V(b0)+2 V(cin)+4 V(a1)+6 V(b1)+8 V(c2)+10
plot V(a0) V(b0)+2 V(cin)+4 V(a1)+6 V(b1)+8 V(a_374_87#)+10

.endc
.end