magic
tech scmos
timestamp 1733169640
<< nwell >>
rect -193 62 -48 115
rect -35 62 -10 115
rect 4 62 29 115
rect 48 41 72 93
<< ntransistor >>
rect 59 10 61 30
rect -182 -11 -180 9
rect -170 -11 -168 9
rect -158 -11 -156 9
rect -146 -11 -144 9
rect -134 -11 -132 9
rect -122 -11 -120 9
rect -110 -11 -108 9
rect -98 -11 -96 9
rect -86 -11 -84 9
rect -74 -11 -72 9
rect -62 -11 -60 9
rect -24 -11 -22 9
rect 15 -11 17 9
<< ptransistor >>
rect -182 68 -180 108
rect -170 68 -168 108
rect -158 68 -156 108
rect -146 68 -144 108
rect -134 68 -132 108
rect -122 68 -120 108
rect -110 68 -108 108
rect -98 68 -96 108
rect -86 68 -84 108
rect -74 68 -72 108
rect -62 68 -60 108
rect -24 68 -22 108
rect 15 68 17 108
rect 59 47 61 87
<< ndiffusion >>
rect 58 10 59 30
rect 61 10 62 30
rect -183 -11 -182 9
rect -180 -11 -179 9
rect -171 -11 -170 9
rect -168 -11 -167 9
rect -159 -11 -158 9
rect -156 -11 -155 9
rect -147 -11 -146 9
rect -144 -11 -143 9
rect -135 -11 -134 9
rect -132 -11 -131 9
rect -123 -11 -122 9
rect -120 -11 -119 9
rect -111 -11 -110 9
rect -108 -11 -107 9
rect -99 -11 -98 9
rect -96 -11 -95 9
rect -87 -11 -86 9
rect -84 -11 -83 9
rect -75 -11 -74 9
rect -72 -11 -71 9
rect -63 -11 -62 9
rect -60 -11 -59 9
rect -25 -11 -24 9
rect -22 -11 -21 9
rect 14 -11 15 9
rect 17 -11 18 9
<< pdiffusion >>
rect -183 68 -182 108
rect -180 68 -179 108
rect -171 68 -170 108
rect -168 68 -167 108
rect -159 68 -158 108
rect -156 68 -155 108
rect -147 68 -146 108
rect -144 68 -143 108
rect -135 68 -134 108
rect -132 68 -131 108
rect -123 68 -122 108
rect -120 68 -119 108
rect -111 68 -110 108
rect -108 68 -107 108
rect -99 68 -98 108
rect -96 68 -95 108
rect -87 68 -86 108
rect -84 68 -83 108
rect -75 68 -74 108
rect -72 68 -71 108
rect -63 68 -62 108
rect -60 68 -59 108
rect -25 68 -24 108
rect -22 68 -21 108
rect 14 68 15 108
rect 17 68 18 108
rect 58 47 59 87
rect 61 47 62 87
<< ndcontact >>
rect 54 10 58 30
rect 62 10 66 30
rect -187 -11 -183 9
rect -179 -11 -171 9
rect -167 -11 -159 9
rect -155 -11 -147 9
rect -143 -11 -135 9
rect -131 -11 -123 9
rect -119 -11 -111 9
rect -107 -11 -99 9
rect -95 -11 -87 9
rect -83 -11 -75 9
rect -71 -11 -63 9
rect -59 -11 -55 9
rect -29 -11 -25 9
rect -21 -11 -17 9
rect 10 -11 14 9
rect 18 -11 22 9
<< pdcontact >>
rect -187 68 -183 108
rect -179 68 -171 108
rect -167 68 -159 108
rect -155 68 -147 108
rect -143 68 -135 108
rect -131 68 -123 108
rect -119 68 -111 108
rect -107 68 -99 108
rect -95 68 -87 108
rect -83 68 -75 108
rect -71 68 -63 108
rect -59 68 -55 108
rect -29 68 -25 108
rect -21 68 -17 108
rect 10 68 14 108
rect 18 68 22 108
rect 54 47 58 87
rect 62 47 66 87
<< polysilicon >>
rect -182 108 -180 111
rect -170 108 -168 111
rect -158 108 -156 111
rect -146 108 -144 111
rect -134 108 -132 111
rect -122 108 -120 111
rect -110 108 -108 111
rect -98 108 -96 111
rect -86 108 -84 111
rect -74 108 -72 111
rect -62 108 -60 111
rect -24 108 -22 111
rect 15 108 17 111
rect 59 87 61 93
rect -182 9 -180 68
rect -170 9 -168 68
rect -158 9 -156 68
rect -146 9 -144 68
rect -134 9 -132 68
rect -122 9 -120 68
rect -110 9 -108 68
rect -98 9 -96 68
rect -86 9 -84 68
rect -74 9 -72 68
rect -62 9 -60 68
rect -24 9 -22 68
rect 15 9 17 68
rect 59 30 61 47
rect 59 6 61 10
rect -182 -16 -180 -11
rect -170 -16 -168 -11
rect -158 -16 -156 -11
rect -146 -15 -144 -11
rect -134 -15 -132 -11
rect -122 -16 -120 -11
rect -110 -16 -108 -11
rect -98 -16 -96 -11
rect -86 -15 -84 -11
rect -74 -15 -72 -11
rect -62 -15 -60 -11
rect -24 -15 -22 -11
rect 15 -15 17 -11
<< polycontact >>
rect 54 34 59 38
<< metal1 >>
rect -193 115 72 119
rect -28 60 -25 68
rect -21 60 -17 68
rect 11 60 14 68
rect 18 60 22 68
rect 54 87 57 115
rect 62 38 66 47
rect 40 34 54 38
rect 62 34 79 38
rect 62 30 66 34
rect 54 -28 58 10
rect -187 -33 72 -28
<< labels >>
rlabel metal1 59 -30 59 -30 1 gnd
rlabel metal1 59 118 59 118 5 vdd
<< end >>
