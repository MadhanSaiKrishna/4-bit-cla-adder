magic
tech scmos
timestamp 1732015684
<< nwell >>
rect -6 32 18 65
<< ntransistor >>
rect 5 0 7 10
<< ptransistor >>
rect 5 38 7 58
<< ndiffusion >>
rect 4 0 5 10
rect 7 0 8 10
<< pdiffusion >>
rect 4 38 5 58
rect 7 38 8 58
<< ndcontact >>
rect 0 0 4 10
rect 8 0 12 10
<< pdcontact >>
rect 0 38 4 58
rect 8 38 12 58
<< polysilicon >>
rect 5 58 7 61
rect 5 10 7 38
rect 5 -3 7 0
<< polycontact >>
rect -1 18 5 23
<< metal1 >>
rect 0 61 12 65
rect 0 58 4 61
rect 8 23 12 38
rect -7 18 -1 23
rect 8 18 18 23
rect 8 10 12 18
rect 0 -3 4 0
rect 0 -7 12 -3
<< labels >>
rlabel metal1 6 64 6 64 5 vdd
rlabel metal1 7 -5 7 -5 1 gnd
rlabel metal1 -5 20 -5 20 3 in
rlabel metal1 15 21 15 21 7 out
<< end >>
