magic
tech scmos
timestamp 1733233777
<< nwell >>
rect 316 57 424 109
rect 441 57 465 109
rect 526 40 550 92
<< ntransistor >>
rect 537 9 539 29
rect 327 -75 329 -55
rect 339 -75 341 -55
rect 351 -75 353 -55
rect 363 -75 365 -55
rect 375 -75 377 -55
rect 387 -75 389 -55
rect 399 -75 401 -55
rect 411 -75 413 -55
rect 452 -75 454 -55
<< ptransistor >>
rect 327 63 329 103
rect 339 63 341 103
rect 351 63 353 103
rect 363 63 365 103
rect 375 63 377 103
rect 387 63 389 103
rect 399 63 401 103
rect 411 63 413 103
rect 452 63 454 103
rect 537 46 539 86
<< ndiffusion >>
rect 536 9 537 29
rect 539 9 540 29
rect 326 -75 327 -55
rect 329 -75 330 -55
rect 338 -75 339 -55
rect 341 -75 342 -55
rect 350 -75 351 -55
rect 353 -75 354 -55
rect 362 -75 363 -55
rect 365 -75 366 -55
rect 374 -75 375 -55
rect 377 -75 378 -55
rect 386 -75 387 -55
rect 389 -75 390 -55
rect 398 -75 399 -55
rect 401 -75 402 -55
rect 410 -75 411 -55
rect 413 -75 414 -55
rect 451 -75 452 -55
rect 454 -75 455 -55
<< pdiffusion >>
rect 326 63 327 103
rect 329 63 330 103
rect 338 63 339 103
rect 341 63 342 103
rect 350 63 351 103
rect 353 63 354 103
rect 362 63 363 103
rect 365 63 366 103
rect 374 63 375 103
rect 377 63 378 103
rect 386 63 387 103
rect 389 63 390 103
rect 398 63 399 103
rect 401 63 402 103
rect 410 63 411 103
rect 413 63 414 103
rect 451 63 452 103
rect 454 63 455 103
rect 536 46 537 86
rect 539 46 540 86
<< ndcontact >>
rect 532 9 536 29
rect 540 9 544 29
rect 322 -75 326 -55
rect 330 -75 338 -55
rect 342 -75 350 -55
rect 354 -75 362 -55
rect 366 -75 374 -55
rect 378 -75 386 -55
rect 390 -75 398 -55
rect 402 -75 410 -55
rect 414 -75 418 -55
rect 447 -75 451 -55
rect 455 -75 459 -55
<< pdcontact >>
rect 322 63 326 103
rect 330 63 338 103
rect 342 63 350 103
rect 354 63 362 103
rect 366 63 374 103
rect 378 63 386 103
rect 390 63 398 103
rect 402 63 410 103
rect 414 63 418 103
rect 447 63 451 103
rect 455 63 459 103
rect 532 46 536 86
rect 540 46 544 86
<< polysilicon >>
rect 327 103 329 106
rect 339 103 341 106
rect 351 103 353 106
rect 363 103 365 106
rect 375 103 377 106
rect 387 103 389 106
rect 399 103 401 106
rect 411 103 413 106
rect 452 103 454 107
rect 537 86 539 92
rect 327 -55 329 63
rect 339 -55 341 63
rect 351 -55 353 63
rect 363 -55 365 63
rect 375 -55 377 63
rect 387 -55 389 63
rect 399 -55 401 63
rect 411 -55 413 63
rect 452 -55 454 63
rect 537 29 539 46
rect 537 5 539 9
rect 327 -79 329 -75
rect 339 -79 341 -75
rect 351 -79 353 -75
rect 363 -79 365 -75
rect 375 -79 377 -75
rect 387 -79 389 -75
rect 399 -79 401 -75
rect 411 -79 413 -75
rect 452 -79 454 -75
<< polycontact >>
rect 323 25 327 29
rect 335 16 339 20
rect 353 8 358 12
rect 358 0 363 4
rect 371 -9 375 -5
rect 383 -17 387 -13
rect 395 -26 399 -22
rect 407 -33 411 -29
rect 532 33 537 37
<< metal1 >>
rect 322 120 535 124
rect 322 103 326 120
rect 381 103 385 120
rect 392 111 451 115
rect 392 103 396 111
rect 447 103 451 111
rect 344 39 347 63
rect 356 54 360 63
rect 404 55 408 63
rect 356 50 403 54
rect 414 37 418 63
rect 455 55 459 63
rect 532 86 535 120
rect 540 37 544 46
rect 349 34 532 37
rect 306 25 316 29
rect 321 25 323 29
rect 306 16 335 20
rect 323 12 327 16
rect 323 8 353 12
rect 308 0 358 4
rect 308 -9 356 -5
rect 361 -9 371 -5
rect 308 -17 383 -13
rect 361 -26 395 -22
rect 321 -33 407 -29
rect 344 -55 347 -47
rect 356 -49 403 -45
rect 356 -55 360 -49
rect 404 -55 408 -49
rect 414 -55 418 34
rect 540 33 560 37
rect 540 29 544 33
rect 435 -49 459 -45
rect 455 -55 459 -49
rect 322 -86 326 -75
rect 380 -86 384 -75
rect 393 -80 396 -75
rect 447 -80 451 -75
rect 393 -83 451 -80
rect 532 -86 536 9
rect 322 -91 536 -86
<< m2contact >>
rect 403 50 408 55
rect 343 34 349 39
rect 455 50 460 55
rect 316 24 321 30
rect 356 -9 361 -4
rect 356 -26 361 -21
rect 315 -33 321 -28
rect 343 -47 348 -42
rect 403 -49 409 -44
rect 428 -49 435 -44
<< metal2 >>
rect 408 50 455 54
rect 316 -28 320 24
rect 344 -42 347 34
rect 356 -21 360 -9
rect 409 -49 428 -45
rect 435 -49 436 -45
<< labels >>
rlabel metal1 510 120 519 124 5 vdd
rlabel metal1 548 33 553 37 1 c2
rlabel metal1 489 -90 496 -87 1 gnd
rlabel metal1 315 26 318 29 3 a1
rlabel metal1 316 16 320 20 3 b1
rlabel metal1 317 0 320 4 3 b0
rlabel metal1 317 -9 320 -5 3 a0
rlabel metal1 317 -17 320 -13 3 cin
<< end >>
