magic
tech scmos
timestamp 1733286918
<< nwell >>
rect 222 151 246 203
rect 266 111 326 203
rect 385 112 409 164
rect 183 44 207 96
rect 429 72 489 164
rect 497 85 534 184
rect 547 87 573 184
rect 593 87 619 184
rect 625 88 653 140
rect 346 5 370 57
<< ntransistor >>
rect 233 120 235 140
rect 396 81 398 101
rect 194 13 196 33
rect 277 12 279 52
rect 289 12 291 52
rect 301 12 303 52
rect 313 12 315 52
rect 640 57 642 77
rect 357 -26 359 -6
rect 440 -27 442 13
rect 452 -27 454 13
rect 464 -27 466 13
rect 476 -27 478 13
rect 509 9 511 49
rect 560 12 562 52
rect 572 12 574 52
rect 606 12 608 52
rect 618 12 620 52
<< ptransistor >>
rect 233 157 235 197
rect 277 117 279 197
rect 289 117 291 197
rect 301 117 303 197
rect 313 117 315 197
rect 396 118 398 158
rect 194 50 196 90
rect 440 78 442 158
rect 452 78 454 158
rect 464 78 466 158
rect 476 78 478 158
rect 509 93 511 173
rect 521 93 523 173
rect 560 93 562 173
rect 606 93 608 173
rect 640 94 642 134
rect 357 11 359 51
<< ndiffusion >>
rect 232 120 233 140
rect 235 120 236 140
rect 395 81 396 101
rect 398 81 399 101
rect 193 13 194 33
rect 196 13 197 33
rect 276 12 277 52
rect 279 12 280 52
rect 288 12 289 52
rect 291 12 292 52
rect 300 12 301 52
rect 303 14 304 52
rect 312 14 313 52
rect 303 12 313 14
rect 315 12 316 52
rect 639 57 640 77
rect 642 57 643 77
rect 356 -26 357 -6
rect 359 -26 360 -6
rect 439 -27 440 13
rect 442 -27 443 13
rect 451 -27 452 13
rect 454 -27 455 13
rect 463 -27 464 13
rect 466 -25 467 13
rect 475 -25 476 13
rect 466 -27 476 -25
rect 478 -27 479 13
rect 508 9 509 49
rect 511 9 512 49
rect 559 12 560 52
rect 562 12 563 52
rect 571 12 572 52
rect 574 12 575 52
rect 605 12 606 52
rect 608 12 609 52
rect 617 12 618 52
rect 620 12 621 52
<< pdiffusion >>
rect 232 157 233 197
rect 235 157 236 197
rect 276 117 277 197
rect 279 117 280 197
rect 288 117 289 197
rect 291 117 292 197
rect 300 117 301 197
rect 303 117 304 197
rect 312 117 313 197
rect 315 117 316 197
rect 395 118 396 158
rect 398 118 399 158
rect 193 50 194 90
rect 196 50 197 90
rect 439 78 440 158
rect 442 78 443 158
rect 451 78 452 158
rect 454 78 455 158
rect 463 78 464 158
rect 466 78 467 158
rect 475 78 476 158
rect 478 78 479 158
rect 508 93 509 173
rect 511 93 512 173
rect 520 93 521 173
rect 523 93 524 173
rect 559 93 560 173
rect 562 93 563 173
rect 605 93 606 173
rect 608 93 609 173
rect 639 94 640 134
rect 642 94 643 134
rect 356 11 357 51
rect 359 11 360 51
<< ndcontact >>
rect 228 120 232 140
rect 236 120 240 140
rect 391 81 395 101
rect 399 81 403 101
rect 189 13 193 33
rect 197 13 201 33
rect 272 12 276 52
rect 280 12 288 52
rect 292 12 300 52
rect 304 14 312 52
rect 316 12 320 52
rect 635 57 639 77
rect 643 57 647 77
rect 352 -26 356 -6
rect 360 -26 364 -6
rect 435 -27 439 13
rect 443 -27 451 13
rect 455 -27 463 13
rect 467 -25 475 13
rect 479 -27 483 13
rect 504 9 508 49
rect 512 9 516 49
rect 555 12 559 52
rect 563 12 571 52
rect 575 12 579 52
rect 601 12 605 52
rect 609 12 617 52
rect 621 12 625 52
<< pdcontact >>
rect 228 157 232 197
rect 236 157 240 197
rect 272 117 276 197
rect 280 117 288 197
rect 292 117 300 197
rect 304 117 312 197
rect 316 117 320 197
rect 391 118 395 158
rect 399 118 403 158
rect 189 50 193 90
rect 197 50 201 90
rect 435 78 439 158
rect 443 78 451 158
rect 455 78 463 158
rect 467 78 475 158
rect 479 78 483 158
rect 504 93 508 173
rect 512 93 520 173
rect 524 93 528 173
rect 555 93 559 173
rect 563 93 567 173
rect 601 93 605 173
rect 609 93 613 173
rect 635 94 639 134
rect 643 94 647 134
rect 352 11 356 51
rect 360 11 364 51
<< polysilicon >>
rect 233 197 235 203
rect 277 197 279 201
rect 289 197 291 201
rect 301 197 303 201
rect 313 197 315 201
rect 233 140 235 157
rect 233 116 235 120
rect 509 173 511 177
rect 521 173 523 177
rect 560 173 562 177
rect 606 173 608 177
rect 396 158 398 164
rect 440 158 442 162
rect 452 158 454 162
rect 464 158 466 162
rect 476 158 478 162
rect 194 90 196 96
rect 277 52 279 117
rect 289 52 291 117
rect 301 52 303 117
rect 313 52 315 117
rect 396 101 398 118
rect 396 77 398 81
rect 640 134 642 140
rect 194 33 196 50
rect 194 9 196 13
rect 357 51 359 57
rect 277 8 279 12
rect 289 8 291 12
rect 301 7 303 12
rect 313 7 315 12
rect 440 13 442 78
rect 452 13 454 78
rect 464 13 466 78
rect 476 13 478 78
rect 509 49 511 93
rect 521 69 523 93
rect 560 76 562 93
rect 606 76 608 93
rect 640 77 642 94
rect 560 52 562 63
rect 572 52 574 64
rect 606 52 608 63
rect 618 52 620 64
rect 640 53 642 57
rect 357 -6 359 11
rect 357 -30 359 -26
rect 509 3 511 9
rect 560 8 562 12
rect 572 9 574 12
rect 606 8 608 12
rect 618 9 620 12
rect 440 -31 442 -27
rect 452 -31 454 -27
rect 464 -32 466 -27
rect 476 -32 478 -27
<< polycontact >>
rect 228 144 233 148
rect 271 94 277 98
rect 284 86 289 90
rect 296 76 301 80
rect 309 66 313 70
rect 391 105 396 109
rect 189 37 194 41
rect 434 55 440 59
rect 447 47 452 51
rect 459 37 464 41
rect 472 27 476 31
rect 503 64 509 69
rect 635 80 640 84
rect 523 72 529 76
rect 558 72 564 76
rect 604 72 610 76
rect 559 63 563 67
rect 571 64 575 69
rect 605 63 609 67
rect 617 64 621 69
rect 352 -2 357 2
<< metal1 >>
rect 189 203 326 207
rect 171 144 181 148
rect 189 90 193 203
rect 228 197 232 203
rect 292 197 300 203
rect 236 148 240 157
rect 207 144 228 148
rect 236 144 251 148
rect 208 82 213 144
rect 236 140 240 144
rect 173 37 177 41
rect 197 41 201 50
rect 182 37 189 41
rect 197 37 216 41
rect 197 33 201 37
rect 189 5 193 13
rect 228 5 232 120
rect 247 98 251 144
rect 497 179 639 187
rect 504 173 508 179
rect 555 173 559 179
rect 601 173 605 179
rect 272 109 276 117
rect 316 109 320 117
rect 352 164 489 168
rect 272 105 344 109
rect 272 104 336 105
rect 247 94 271 98
rect 255 86 284 90
rect 254 76 296 80
rect 247 66 309 70
rect 247 42 252 66
rect 272 56 320 61
rect 272 52 276 56
rect 316 52 320 56
rect 304 12 312 14
rect 282 5 286 12
rect 189 1 286 5
rect 306 5 310 12
rect 324 5 328 104
rect 352 51 356 164
rect 391 158 395 164
rect 455 158 463 164
rect 399 109 403 118
rect 370 105 391 109
rect 399 105 414 109
rect 371 43 376 105
rect 399 101 403 105
rect 306 1 328 5
rect 336 -2 340 2
rect 360 2 364 11
rect 345 -2 352 2
rect 360 -2 379 2
rect 360 -6 364 -2
rect 352 -34 356 -26
rect 391 -34 395 81
rect 410 59 414 105
rect 635 134 639 179
rect 524 83 528 93
rect 435 70 439 78
rect 479 70 483 78
rect 512 79 528 83
rect 563 84 567 93
rect 550 80 588 84
rect 609 84 613 93
rect 643 85 647 94
rect 596 80 635 84
rect 643 81 661 85
rect 435 69 499 70
rect 435 65 503 69
rect 410 55 434 59
rect 418 47 447 51
rect 417 37 459 41
rect 410 27 472 31
rect 410 3 415 27
rect 435 17 483 22
rect 435 13 439 17
rect 479 13 483 17
rect 467 -27 475 -25
rect 445 -34 449 -27
rect 352 -38 449 -34
rect 469 -34 473 -27
rect 487 -34 491 65
rect 498 64 503 65
rect 512 67 516 79
rect 529 72 535 76
rect 585 76 588 80
rect 643 77 647 81
rect 540 72 558 76
rect 564 72 582 76
rect 585 72 604 76
rect 610 72 621 76
rect 571 69 575 72
rect 512 63 559 67
rect 578 67 582 72
rect 617 69 621 72
rect 578 63 605 67
rect 512 49 516 63
rect 504 3 508 9
rect 575 3 579 12
rect 621 3 625 12
rect 635 3 640 57
rect 500 -2 640 3
rect 469 -38 491 -34
<< m2contact >>
rect 181 143 186 149
rect 202 144 207 149
rect 208 75 214 82
rect 177 37 182 42
rect 216 36 222 42
rect 344 104 349 110
rect 249 85 255 91
rect 248 74 254 81
rect 246 37 252 42
rect 365 105 370 110
rect 371 36 377 43
rect 340 -2 345 3
rect 379 -3 385 3
rect 545 80 550 85
rect 591 80 596 85
rect 412 46 418 52
rect 411 35 417 42
rect 409 -2 415 3
rect 535 72 540 77
rect 554 52 559 57
rect 600 52 605 57
<< metal2 >>
rect 186 144 202 148
rect 349 105 365 109
rect 178 86 249 90
rect 178 42 182 86
rect 214 76 248 80
rect 535 58 540 72
rect 498 54 540 58
rect 545 57 550 80
rect 591 57 596 80
rect 545 52 554 57
rect 591 52 600 57
rect 341 47 412 51
rect 222 37 246 41
rect 341 3 345 47
rect 377 37 411 41
rect 385 -2 409 2
<< labels >>
rlabel metal1 194 3 194 3 1 gnd
rlabel metal1 194 205 194 205 5 vdd
rlabel metal1 235 3 235 3 1 gnd
rlabel metal1 233 206 233 206 5 vdd
rlabel space 183 36 189 41 1 a0
rlabel metal1 216 144 223 148 1 b0
rlabel space 174 144 181 150 1 b0
rlabel metal1 357 -36 357 -36 1 gnd
rlabel metal1 357 166 357 166 5 vdd
rlabel metal1 398 -36 398 -36 1 gnd
rlabel metal1 396 167 396 167 5 vdd
rlabel metal1 346 -2 351 2 1 c0
rlabel metal1 532 74 532 74 1 clk
rlabel metal1 512 -1 512 -1 1 gnd
rlabel metal1 605 184 605 184 5 vdd
rlabel metal1 559 184 559 184 5 vdd
rlabel metal1 516 185 516 185 5 vdd
rlabel metal2 505 56 505 56 1 clk
rlabel metal1 653 81 658 85 1 s0
rlabel space 493 63 502 71 1 s0_out
<< end >>
