* SPICE3 file created from carry_one.ext - technology: scmos
.include TSMC_180nm.txt
.option scale=0.09u
.param SUPPLY = 1.8
.param LAMBDA=0.09u
.global gnd vdd
Vdd vdd gnd 'SUPPLY'

V1 A0_in gnd pulse 0 1.8 0u 10p 10p 0.1u 0.3u
V2 B0_in gnd pulse 0 1.8 0.3u 10p 10p 0.1u 0.3u
V3 A1_in gnd pulse 0 1.8 0.5u 10p 10p 0.01u 0.03u
V4 B1_in gnd pulse 0 1.8 0u 10p 10p 0.02u 0.03u
V5 A2_in gnd pulse 0 1.8 0.5u 10p 10p 0.1u 0.3u
V6 B2_in gnd pulse 0 1.8 0u 10p 10p 0.1u 0.3u
V7 A3_in gnd pulse 0 1.8 0.5u 10p 10p 0.01u 0.03u
V8 B3_in gnd pulse 0 1.8 0u 10p 10p 0.02u 0.07u

V9 clk gnd pulse 0 1.8 0.03u 10p 10p 60n 100n


V10 Cin gnd dc 0

M1000 a_n7_12# a1_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=12200 ps=4860
M1001 a_1344_n270# a_1300_n267# a_1337_n270# w_1331_n276# CMOSP w=80 l=2
+  ad=800 pd=180 as=800 ps=340
M1002 gnd clk a_374_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1003 a_759_164# a0 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1004 a_1472_n267# cin vdd w_1459_n236# CMOSP w=40 l=2
+  ad=200 pd=90 as=24400 ps=8900
M1005 a_723_455# b2 a_711_164# w_686_449# CMOSP w=40 l=2
+  ad=1000 pd=290 as=600 ps=190
M1006 a_1472_n267# cin gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1007 a_817_889# b0 a_853_889# w_902_883# CMOSP w=40 l=2
+  ad=1000 pd=290 as=600 ps=190
M1008 a_760_37# cin vdd w_687_31# CMOSP w=40 l=2
+  ad=600 pd=190 as=0 ps=0
M1009 a_n125_n236# a_n176_n239# a_n132_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1010 a_712_n101# b1 a_700_n101# Gnd CMOSN w=20 l=2
+  ad=300 pd=110 as=200 ps=60
M1011 vdd a3 a_1354_614# w_1341_608# CMOSP w=80 l=2
+  ad=0 pd=0 as=800 ps=180
M1012 a_1305_329# a2 vdd w_1292_360# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1013 a_1347_37# a_1303_40# a_1340_37# w_1334_31# CMOSP w=80 l=2
+  ad=800 pd=180 as=800 ps=340
M1014 a_1266_222# b2 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1015 n010 a0 a_714_n308# w_677_n314# CMOSP w=40 l=2
+  ad=600 pd=270 as=600 ps=190
M1016 a_1349_326# a_1305_329# a_1342_326# w_1336_320# CMOSP w=80 l=2
+  ad=800 pd=180 as=800 ps=340
M1017 a_699_164# a2 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1018 a1 a_83_15# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1019 a_1538_509# a_1347_614# gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1020 a_721_551# a3 a_733_889# w_941_883# CMOSP w=40 l=2
+  ad=600 pd=190 as=1000 ps=290
M1021 a_724_37# a0 a_760_37# w_687_31# CMOSP w=40 l=2
+  ad=1000 pd=290 as=0 ps=0
M1022 s1_out c1 a_1531_n68# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=400 ps=100
M1023 a_159_96# a_151_67# vdd w_145_88# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1024 vdd a_1337_n270# a_1516_n270# w_1503_n276# CMOSP w=80 l=2
+  ad=0 pd=0 as=800 ps=180
M1025 a_159_12# a_151_67# gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1026 a_1303_40# a1 vdd w_1290_71# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1027 a_255_n236# clk a_248_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1028 a_1550_614# c3 vdd w_1513_608# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1029 a_37_15# clk vdd w_29_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1030 vdd a0 a_829_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1031 a_1361_221# b2 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1032 a_n85_15# a_n131_15# vdd w_n93_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1033 gnd a_n131_15# a_n78_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1034 a_209_n236# a_158_n239# a_202_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1035 vdd b1 a_1347_37# w_1334_31# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 a_n86_n236# a_n132_n236# vdd w_n94_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1037 a_82_n236# a_36_n236# vdd w_74_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1038 vdd a0 a_1344_n270# w_1331_n276# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 cout a_721_551# vdd w_985_824# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1040 a_1366_509# a3 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1041 a_83_15# a_37_15# vdd w_75_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1042 s0_out a_1433_n374# a_1540_n270# w_1503_n276# CMOSP w=80 l=2
+  ad=800 pd=340 as=800 ps=180
M1043 a_1436_n67# a_1340_37# vdd w_1423_n36# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1044 a_781_889# b1 a_769_889# w_692_883# CMOSP w=40 l=2
+  ad=1000 pd=290 as=400 ps=100
M1045 a3 a_414_15# vdd w_438_91# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1046 a_1436_n67# a_1340_37# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1047 a_1271_510# a3 vdd w_1258_541# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1048 a_1477_329# c2 vdd w_1464_360# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1049 a_712_n101# a1 a_724_37# w_687_31# CMOSP w=40 l=2
+  ad=600 pd=190 as=0 ps=0
M1050 a_724_n101# b1 a_712_n101# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=0 ps=0
M1051 a_771_164# b0 a_759_164# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=0 ps=0
M1052 a_735_455# b1 a_723_455# w_686_449# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1053 a_159_12# clk a_159_96# w_145_88# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1054 a_1310_617# b3 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1055 a_723_455# b1 a_771_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=1000 ps=290
M1056 a_44_15# a_n7_12# a_37_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1057 a_n8_n155# b1_in vdd w_n22_n163# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1058 a_1378_614# b3 vdd w_1341_608# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1059 a_733_551# b3 a_721_551# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=300 ps=110
M1060 gnd a_37_15# a_90_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1061 c3 a_711_164# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1062 a_n78_15# clk a_n85_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1063 vdd b2 a_1349_326# w_1336_320# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 a_1371_37# a1 vdd w_1334_31# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1065 a_n8_n239# clk a_n8_n155# w_n22_n163# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1066 b1 a_82_n236# vdd w_106_n160# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1067 a_367_n236# clk vdd w_359_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1068 s3_out c3 a_1538_509# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1069 a_203_15# clk vdd w_195_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1070 a_1433_n374# a_1337_n270# vdd w_1420_n343# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1071 b1 a_82_n236# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1072 a_249_15# a_203_15# vdd w_241_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1073 a_90_15# clk a_83_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1074 a_1433_n374# a_1337_n270# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1075 a_1540_n270# cin vdd w_1503_n276# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 a_1264_n67# b1 vdd w_1251_n36# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1077 a_368_15# clk vdd w_360_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1078 a_1264_n67# b1 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1079 a0 a_n85_15# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1080 a_771_164# b0 a_807_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=300 ps=110
M1081 gnd a_202_n236# a_255_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 a_1512_n68# a_1436_n67# s1_out Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1083 a_1533_221# a_1342_326# gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1084 a2 a_249_15# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1085 gnd clk a_209_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 a_700_37# a1 vdd w_687_31# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1087 a_1340_37# a_1264_n67# a_1371_37# w_1334_31# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 a_1368_n270# b0 vdd w_1331_n276# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1089 a_1300_n267# b0 vdd w_1287_n236# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1090 gnd clk a_44_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 a_1300_n267# b0 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1092 gnd a_367_n236# a_420_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1093 a_711_164# a2 a_723_164# Gnd CMOSN w=20 l=2
+  ad=300 pd=110 as=500 ps=170
M1094 a_690_n370# b0 n010 Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=300 ps=150
M1095 a_736_n101# b0 a_724_n101# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1096 a_1443_510# a_1347_614# vdd w_1430_541# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1097 a_807_455# a0 a_771_455# w_686_449# CMOSP w=40 l=2
+  ad=600 pd=190 as=0 ps=0
M1098 a_210_15# a_159_12# a_203_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1099 a_1347_614# b3 a_1366_509# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1100 a_256_15# clk a_249_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1101 a_781_551# a2 a_733_551# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=0 ps=0
M1102 a_n175_12# clk a_n175_96# w_n189_88# CMOSP w=80 l=2
+  ad=400 pd=170 as=800 ps=180
M1103 a_324_96# a3_in vdd w_310_88# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1104 a_375_15# a_324_12# a_368_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1105 a_1340_n68# a_1264_n67# a_1340_37# Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=400 ps=100
M1106 a_1475_40# c1 vdd w_1462_71# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1107 a_853_551# cin gnd Gnd CMOSN w=20 l=2
+  ad=300 pd=110 as=0 ps=0
M1108 a_324_12# a3_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1109 a_158_n239# b2_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1110 vdd a1 a_735_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 vdd a_1342_326# a_1521_326# w_1508_320# CMOSP w=80 l=2
+  ad=0 pd=0 as=800 ps=180
M1112 a_1347_614# a_1271_510# a_1378_614# w_1341_608# CMOSP w=80 l=2
+  ad=800 pd=340 as=0 ps=0
M1113 a_771_455# a1 a_723_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 gnd clk a_210_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 a_420_n236# clk a_413_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1116 a_733_889# b3 a_721_551# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1117 a_745_551# b2 a_733_551# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1118 a_733_551# b2 a_781_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 a_n132_n236# clk vdd w_n140_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1120 a_323_n239# b3_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1121 a_723_164# b2 a_711_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gnd a_203_15# a_256_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 gnd a_1472_n267# a_1509_n375# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1124 gnd a_1475_40# a_1512_n68# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 s2_out c2 a_1533_221# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1126 a_n175_96# a0_in vdd w_n189_88# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 a_324_12# clk a_324_96# w_310_88# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1128 gnd clk a_375_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 a_1337_n270# a_1261_n374# a_1368_n270# w_1331_n276# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 a_690_n308# b0 n010 w_677_n314# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1131 a_n175_12# a0_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1132 gnd a_1300_n267# a_1337_n375# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1133 gnd a0 a_736_n101# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 a_1303_40# a1 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1135 a_43_n236# a_n8_n239# a_36_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1136 a_248_n236# a_202_n236# vdd w_240_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1137 vdd cin a_807_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 a_202_n236# clk vdd w_194_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1139 a_1347_509# a_1271_510# a_1347_614# Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1140 a_1438_222# a_1342_326# vdd w_1425_253# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1141 gnd a_1303_40# a_1340_n68# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 a_781_889# a2 a_733_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 a_817_551# b1 a_781_551# Gnd CMOSN w=20 l=2
+  ad=500 pd=170 as=0 ps=0
M1144 a_1261_n374# a0 vdd w_1248_n343# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1145 a_1519_37# a_1475_40# s1_out w_1506_31# CMOSP w=80 l=2
+  ad=800 pd=180 as=800 ps=340
M1146 a_711_164# b2 a_699_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1147 gnd clk a_n124_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1148 a_1261_n374# a0 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1149 a_724_n101# a0 a_760_n101# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=300 ps=110
M1150 a_853_889# cin vdd w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 a_1310_617# b3 vdd w_1297_648# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1152 a_817_551# a0 a_853_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 s3_out a_1443_510# a_1550_614# w_1513_608# CMOSP w=80 l=2
+  ad=800 pd=340 as=0 ps=0
M1154 a_1342_326# a2 a_1361_221# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1155 a_n131_15# clk vdd w_n139_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1156 a3 a_414_15# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1157 a_1271_510# a3 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1158 a_759_455# a0 vdd w_686_449# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1159 a_1545_326# c2 vdd w_1508_320# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1160 a_414_15# a_368_15# vdd w_406_90# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1161 gnd a0 a_690_n370# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 a_709_551# a3 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1163 c3 a_711_164# vdd w_919_379# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1164 a_724_37# a_823_n105# a_760_37# w_812_31# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 a_n176_n239# b0_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1166 a_745_889# b2 a_733_889# w_692_883# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1167 gnd a2 a_745_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 a_n7_12# clk a_n7_96# w_n21_88# CMOSP w=80 l=2
+  ad=400 pd=170 as=800 ps=180
M1169 a_1482_617# c3 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1170 a_1528_n375# a_1337_n270# gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1171 a_733_889# b2 a_781_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 a_712_n101# b1 a_700_37# w_687_31# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 a_699_455# a2 vdd w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 a_735_164# b1 a_723_164# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1175 b0 a_n86_n236# vdd w_n62_n160# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1176 b0 a_n86_n236# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1177 a_723_164# b1 a_771_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 a_1531_n68# a_1340_37# gnd Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 a_1266_222# b2 vdd w_1253_253# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1180 a_1356_n375# a0 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1181 a_760_n101# cin gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 vdd a_1340_37# a_1519_37# w_1506_31# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 gnd clk a_43_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1184 a_1305_329# a2 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1185 a_1514_221# a_1438_222# s2_out Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1186 a1 a_83_15# vdd w_107_91# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1187 a_n124_15# a_n175_12# a_n131_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1188 a_421_15# clk a_414_15# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1189 a_1509_n375# a_1433_n374# s0_out Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=100
M1190 a_1373_326# a2 vdd w_1336_320# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1191 a_1519_509# a_1443_510# s3_out Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1192 a_158_n155# b2_in vdd w_144_n163# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1193 a_724_37# b1 a_712_n101# w_687_31# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 c1 n010 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1195 a_712_n101# a1 a_724_n101# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 a_1543_37# c1 vdd w_1506_31# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1197 c2 a_712_n101# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1198 vdd a0 a_690_n308# w_677_n314# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1199 a_1443_510# a_1347_614# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1200 gnd a_368_15# a_421_15# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1201 a_n79_n236# clk a_n86_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1202 a_89_n236# clk a_82_n236# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=200 ps=90
M1203 cout a_721_551# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1204 a_829_551# b0 a_817_551# Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1205 a_1526_614# a_1482_617# s3_out w_1513_608# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1206 a_714_n370# cin gnd Gnd CMOSN w=20 l=2
+  ad=300 pd=110 as=0 ps=0
M1207 a_1359_n68# b1 gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1208 a_817_889# b1 a_781_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 a_323_n155# b3_in vdd w_309_n163# CMOSP w=80 l=2
+  ad=800 pd=180 as=0 ps=0
M1210 a_781_551# a1 a_817_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1211 a_n176_n239# clk a_n176_n155# w_n190_n163# CMOSP w=80 l=2
+  ad=400 pd=170 as=800 ps=180
M1212 a_817_889# a0 a_853_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 a_771_455# b0 a_759_455# w_686_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 a_1342_221# a_1266_222# a_1342_326# Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1215 a_807_164# a0 a_771_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 s0_out cin a_1528_n375# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 a_1475_40# c1 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1218 a_709_889# a3 vdd w_692_883# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1219 a_721_551# b3 a_709_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1220 s2_out a_1438_222# a_1545_326# w_1508_320# CMOSP w=80 l=2
+  ad=800 pd=340 as=0 ps=0
M1221 a_700_n101# a1 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1222 vdd a2 a_745_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 a_769_551# a1 gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1224 a_724_n101# a_823_n105# a_760_n101# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 a_1477_329# c2 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1226 gnd a1 a_735_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 a_413_n236# a_367_n236# vdd w_405_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1228 a_817_551# b0 a_853_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 a_736_37# b0 a_724_37# w_687_31# CMOSP w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1230 a_1337_n270# b0 a_1356_n375# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1231 n010 b0 a_714_n370# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 s1_out a_1436_n67# a_1543_37# w_1506_31# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1233 a_771_164# a1 a_723_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1234 gnd a_n132_n236# a_n79_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 gnd a_1477_329# a_1514_221# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1236 a_374_n236# a_323_n239# a_367_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1237 a_1354_614# a_1310_617# a_1347_614# w_1341_608# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1238 a_771_455# b0 a_807_455# w_844_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 c2 a_712_n101# vdd w_868_14# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1240 gnd a_1482_617# a_1519_509# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1241 gnd clk a_n125_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1242 a_158_n239# clk a_158_n155# w_144_n163# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1243 a_1342_326# a_1266_222# a_1373_326# w_1336_320# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1244 a_721_551# a3 a_733_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1245 a0 a_n85_15# vdd w_n61_91# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1246 a_714_n308# cin vdd w_677_n314# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1247 gnd a_36_n236# a_89_n236# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1248 a_n8_n239# b1_in gnd Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1249 a2 a_249_15# vdd w_273_91# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1250 n010 a0 a_714_n370# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 b2 a_248_n236# vdd w_272_n160# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1252 a_711_164# a2 a_723_455# w_883_449# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1253 a_36_n236# clk vdd w_28_n161# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1254 b2 a_248_n236# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1255 a_n176_n155# b0_in vdd w_n190_n163# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 a_323_n239# clk a_323_n155# w_309_n163# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1257 vdd a0 a_736_37# w_687_31# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 gnd a0 a_829_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 vdd a_1347_614# a_1526_614# w_1513_608# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 a_1340_37# a1 a_1359_n68# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1261 a_829_889# b0 a_817_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1262 gnd a_1305_329# a_1342_221# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 a_1438_222# a_1342_326# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1264 a_1516_n270# a_1472_n267# s0_out w_1503_n276# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 b3 a_413_n236# vdd w_437_n160# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1266 a_1521_326# a_1477_329# s2_out w_1508_320# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 c1 n010 vdd w_782_n313# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1268 b3 a_413_n236# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1269 a_781_889# a1 a_817_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1270 gnd cin a_807_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 a_721_551# b3 a_709_889# w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1272 gnd a_1310_617# a_1347_509# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 n010 b0 a_714_n308# w_749_n314# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1274 a_1482_617# c3 vdd w_1469_648# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1275 a_781_551# b1 a_769_551# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1276 a_n7_96# a1_in vdd w_n21_88# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1277 a_1337_n375# a_1261_n374# a_1337_n270# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1278 a_769_889# a1 vdd w_692_883# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 a_711_164# b2 a_699_164# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 gnd a_1342_221# 0.52fF
C1 b2 a_1305_329# 0.40fF
C2 gnd a_1528_n375# 0.41fF
C3 w_29_90# clk 0.07fF
C4 gnd a1_in 0.02fF
C5 clk a_n132_n236# 0.85fF
C6 b0 w_n62_n160# 0.06fF
C7 vdd w_1462_71# 0.08fF
C8 vdd a_1340_37# 0.14fF
C9 w_1430_541# a_1443_510# 0.06fF
C10 a_1509_n375# a_1528_n375# 0.08fF
C11 vdd a_1349_326# 0.88fF
C12 vdd a_700_37# 0.41fF
C13 a_721_551# cout 0.05fF
C14 b0_in a_n176_n239# 0.07fF
C15 w_1290_71# a_1303_40# 0.06fF
C16 vdd a_1475_40# 0.44fF
C17 a_1514_221# a_1533_221# 0.08fF
C18 b2 a_733_889# 0.15fF
C19 clk a_367_n236# 0.85fF
C20 gnd a_255_n236# 0.41fF
C21 a2 a_721_551# 0.32fF
C22 w_28_n161# clk 0.07fF
C23 a_1443_510# a_1482_617# 0.08fF
C24 vdd w_272_n160# 0.06fF
C25 vdd w_1248_n343# 0.06fF
C26 a_723_455# a_735_455# 0.41fF
C27 a_368_15# vdd 0.86fF
C28 w_310_88# a_324_12# 0.11fF
C29 b0 a_781_889# 0.10fF
C30 a1 a_733_551# 0.21fF
C31 vdd w_868_14# 0.06fF
C32 cin a_1472_n267# 0.13fF
C33 w_1506_31# a_1436_n67# 0.07fF
C34 a_711_164# a_723_164# 0.96fF
C35 a_n132_n236# a_n125_n236# 0.41fF
C36 c2 a_1438_222# 0.56fF
C37 a_1477_329# a_1342_326# 0.40fF
C38 vdd a_736_37# 0.41fF
C39 vdd cout 0.41fF
C40 vdd w_677_n314# 0.03fF
C41 a_1310_617# w_1341_608# 0.07fF
C42 b0 a_1337_n270# 0.09fF
C43 c2 c1 0.25fF
C44 vdd w_195_90# 0.17fF
C45 a2 vdd 1.54fF
C46 gnd a_n79_n236# 0.41fF
C47 b0 w_749_n314# 0.10fF
C48 b1_in a_n8_n239# 0.07fF
C49 a_853_889# w_692_883# 0.03fF
C50 w_n139_90# a_n131_15# 0.10fF
C51 b2 w_1336_320# 0.07fF
C52 a_711_164# w_686_449# 0.03fF
C53 gnd a_1433_n374# 0.33fF
C54 a_1344_n270# w_1331_n276# 0.02fF
C55 a_1303_40# a_1264_n67# 0.08fF
C56 b2 w_692_883# 0.13fF
C57 w_74_n161# a_82_n236# 0.10fF
C58 a_249_15# a_256_15# 0.41fF
C59 a_733_889# a_745_889# 0.41fF
C60 a_1509_n375# a_1433_n374# 0.43fF
C61 a_1347_614# a_1443_510# 0.20fF
C62 a_1368_n270# a_1337_n270# 0.82fF
C63 a_1538_509# gnd 0.41fF
C64 s3_out a_1526_614# 0.82fF
C65 vdd w_194_n161# 0.17fF
C66 vdd a_n176_n155# 0.88fF
C67 a_711_164# b2 0.18fF
C68 a_712_n101# a_700_n101# 0.21fF
C69 gnd a_1436_n67# 0.33fF
C70 a_1264_n67# a_1340_n68# 0.43fF
C71 w_1513_608# a_1550_614# 0.02fF
C72 a_151_67# a_159_12# 0.07fF
C73 a_771_455# b1 0.01fF
C74 b2 c2 0.14fF
C75 a_159_96# a_159_12# 0.82fF
C76 a_723_455# cin 0.08fF
C77 a2 a_1266_222# 0.56fF
C78 b1 a_1340_37# 0.09fF
C79 w_144_n163# a_158_n239# 0.11fF
C80 gnd a_712_n101# 0.04fF
C81 a_724_37# a_736_37# 0.41fF
C82 vdd a_1371_37# 0.88fF
C83 a0 n010 0.01fF
C84 gnd a_759_164# 0.21fF
C85 a_721_551# w_985_824# 0.08fF
C86 a3_in a_324_12# 0.07fF
C87 a_733_889# w_941_883# 0.06fF
C88 a1 a_712_n101# 0.19fF
C89 s0_out vdd 0.05fF
C90 b0 a_723_164# 0.15fF
C91 a_n7_96# a_n7_12# 0.82fF
C92 vdd a_769_889# 0.41fF
C93 vdd a_1354_614# 0.88fF
C94 a_1340_n68# a_1359_n68# 0.08fF
C95 a_n8_n155# a_n8_n239# 0.82fF
C96 a1 a_817_551# 0.12fF
C97 vdd w_1425_253# 0.06fF
C98 a_1347_509# a_1310_617# 0.09fF
C99 s3_out a_1482_617# 0.12fF
C100 b0 c1 0.15fF
C101 w_n140_n161# a_n132_n236# 0.10fF
C102 a_1514_221# a_1477_329# 0.09fF
C103 a_1361_221# a_1342_326# 0.41fF
C104 a_745_889# w_692_883# 0.02fF
C105 b3 w_437_n160# 0.06fF
C106 gnd a_90_15# 0.41fF
C107 gnd a_700_n101# 0.21fF
C108 vdd a_82_n236# 0.86fF
C109 a_420_n236# a_413_n236# 0.41fF
C110 b0 w_686_449# 0.06fF
C111 vdd w_273_91# 0.06fF
C112 s1_out a_1436_n67# 0.09fF
C113 w_1459_n236# a_1472_n267# 0.06fF
C114 w_1331_n276# a_1337_n270# 0.21fF
C115 w_1506_31# s1_out 0.21fF
C116 vdd w_985_824# 0.06fF
C117 vdd w_1290_71# 0.08fF
C118 w_309_n163# clk 0.08fF
C119 a1 gnd 0.74fF
C120 b3 c3 0.14fF
C121 c3 a_1482_617# 0.13fF
C122 a_1337_n270# a_1433_n374# 0.20fF
C123 a2 a_781_551# 0.09fF
C124 gnd a_1509_n375# 0.52fF
C125 w_1508_320# a_1477_329# 0.07fF
C126 a_n175_12# a0_in 0.07fF
C127 a2 b1 2.13fF
C128 b2 b0 1.09fF
C129 b3 a0 0.89fF
C130 b3 a3 1.97fF
C131 w_437_n160# a_413_n236# 0.08fF
C132 a_n7_12# a_37_15# 0.13fF
C133 a0 cin 5.13fF
C134 cin a3 0.47fF
C135 a_1347_614# s3_out 0.09fF
C136 b2 a_1342_221# 0.09fF
C137 a_735_455# vdd 0.41fF
C138 vdd n010 0.39fF
C139 w_1513_608# a_1443_510# 0.07fF
C140 gnd a_43_n236# 0.41fF
C141 vdd a_1342_326# 0.14fF
C142 vdd w_1503_n276# 0.09fF
C143 a_n175_96# w_n189_88# 0.02fF
C144 w_272_n160# a_248_n236# 0.08fF
C145 gnd s1_out 0.15fF
C146 a_714_n308# w_677_n314# 0.03fF
C147 w_28_n161# a_36_n236# 0.10fF
C148 vdd a_1264_n67# 0.41fF
C149 clk a_202_n236# 0.85fF
C150 b3 a_721_551# 0.17fF
C151 a_1347_614# c3 0.57fF
C152 vdd a_1526_614# 0.88fF
C153 a_711_164# a_723_455# 1.40fF
C154 a_368_15# w_360_90# 0.10fF
C155 a_203_15# vdd 0.86fF
C156 cin a_721_551# 0.17fF
C157 a1 a_781_889# 0.10fF
C158 a0 a_733_889# 0.15fF
C159 vdd a_159_12# 0.03fF
C160 vdd w_1287_n236# 0.08fF
C161 b2 a_733_551# 0.21fF
C162 a_1347_614# a3 0.09fF
C163 vdd w_1430_541# 0.06fF
C164 a_n7_12# vdd 0.03fF
C165 w_902_883# b0 0.06fF
C166 gnd a_n125_n236# 0.41fF
C167 c2 a_1477_329# 0.13fF
C168 a_1266_222# a_1342_326# 0.09fF
C169 gnd a_1337_n270# 0.26fF
C170 vdd a_829_889# 0.41fF
C171 b1 a_82_n236# 0.05fF
C172 a_1342_326# s2_out 0.09fF
C173 a_n176_n155# a_n176_n239# 0.82fF
C174 vdd w_107_91# 0.06fF
C175 b3 vdd 1.44fF
C176 vdd a_1482_617# 0.44fF
C177 a_1340_37# a_1475_40# 0.40fF
C178 a_1509_n375# a_1337_n270# 0.09fF
C179 a_1436_n67# c1 0.56fF
C180 w_n189_88# clk 0.08fF
C181 w_1462_71# a_1475_40# 0.06fF
C182 w_1251_n36# a_1264_n67# 0.06fF
C183 w_1506_31# c1 0.07fF
C184 a_1344_n270# a_1337_n270# 0.82fF
C185 a0 w_687_31# 0.13fF
C186 cin vdd 0.84fF
C187 a_203_15# a_210_15# 0.41fF
C188 a_807_455# w_686_449# 0.03fF
C189 a_771_455# w_844_449# 0.06fF
C190 a_1337_n375# a0 0.09fF
C191 a_721_551# a_733_889# 1.48fF
C192 vdd a_1543_37# 0.88fF
C193 a0 w_692_883# 0.13fF
C194 vdd a_1305_329# 0.44fF
C195 a3 w_692_883# 0.06fF
C196 a_1366_509# gnd 0.41fF
C197 a_1436_n67# a_1512_n68# 0.43fF
C198 w_310_88# clk 0.08fF
C199 a_89_n236# a_82_n236# 0.41fF
C200 vdd w_106_n160# 0.06fF
C201 a_711_164# c3 0.05fF
C202 w_1513_608# s3_out 0.21fF
C203 c3 c2 0.26fF
C204 a_711_164# a0 0.26fF
C205 a_723_455# b0 0.15fF
C206 gnd a_1438_222# 0.33fF
C207 gnd a_421_15# 0.41fF
C208 a1 w_1334_31# 0.07fF
C209 vdd a_413_n236# 0.86fF
C210 a0 c2 0.14fF
C211 a_1337_n375# a_1261_n374# 0.43fF
C212 a3 c2 0.14fF
C213 gnd c1 0.44fF
C214 a1 a_723_164# 0.15fF
C215 a_83_15# a_90_15# 0.41fF
C216 a_1354_614# w_1341_608# 0.02fF
C217 vdd a_1347_614# 0.14fF
C218 a_1305_329# a_1266_222# 0.08fF
C219 cin a_724_37# 0.08fF
C220 vdd w_1508_320# 0.09fF
C221 cin a_771_164# 0.01fF
C222 b1 a_1264_n67# 0.20fF
C223 a1 c1 0.15fF
C224 a_721_551# w_692_883# 0.03fF
C225 a3_in gnd 0.02fF
C226 gnd a_249_15# 0.10fF
C227 a0 a_853_551# 0.09fF
C228 w_1513_608# c3 0.07fF
C229 w_1258_541# a_1271_510# 0.06fF
C230 a_n7_12# w_n21_88# 0.11fF
C231 w_241_90# a_249_15# 0.10fF
C232 a_1514_221# s2_out 1.02fF
C233 vdd a_n8_n155# 0.89fF
C234 a_83_15# gnd 0.10fF
C235 gnd a_1512_n68# 0.52fF
C236 a_1472_n267# a_1433_n374# 0.08fF
C237 a1 w_686_449# 0.13fF
C238 a_n85_15# a0 0.05fF
C239 a_83_15# a1 0.05fF
C240 a_1371_37# a_1340_37# 0.82fF
C241 w_240_n161# a_202_n236# 0.07fF
C242 a_714_n308# n010 1.06fF
C243 vdd w_687_31# 0.10fF
C244 w_1287_n236# a_1300_n267# 0.06fF
C245 cin a_724_n101# 0.08fF
C246 b2 gnd 0.96fF
C247 b3 a_1310_617# 0.13fF
C248 a1 a_853_889# 0.09fF
C249 w_n140_n161# clk 0.07fF
C250 vdd w_1336_320# 0.09fF
C251 w_1464_360# c2 0.08fF
C252 b2 a1 1.34fF
C253 a_249_15# clk 0.13fF
C254 vdd a_158_n239# 0.03fF
C255 vdd w_692_883# 0.14fF
C256 b3 b1 0.82fF
C257 s1_out c1 0.09fF
C258 b0 c3 0.14fF
C259 cin a_781_551# 0.09fF
C260 a3 a_1271_510# 0.20fF
C261 w_1508_320# s2_out 0.21fF
C262 a_83_15# clk 0.13fF
C263 b0 a0 7.29fF
C264 b1 cin 0.89fF
C265 a_158_n155# a_158_n239# 0.82fF
C266 vdd w_1459_n236# 0.08fF
C267 b0 a3 1.93fF
C268 gnd a_1533_221# 0.41fF
C269 w_145_88# clk 0.08fF
C270 s1_out a_1512_n68# 1.02fF
C271 w_29_90# a_37_15# 0.10fF
C272 w_782_n313# n010 0.08fF
C273 vdd c2 1.11fF
C274 b1 w_106_n160# 0.06fF
C275 vdd w_1423_n36# 0.06fF
C276 w_1336_320# a_1266_222# 0.07fF
C277 vdd a_1521_326# 0.88fF
C278 w_687_31# a_724_37# 0.06fF
C279 w_n22_n163# b1_in 0.08fF
C280 b0 a_1261_n374# 0.56fF
C281 a_1342_221# a_1361_221# 0.08fF
C282 a_714_n370# gnd 0.21fF
C283 clk a_36_n236# 0.85fF
C284 a_781_889# a_853_889# 0.16fF
C285 a_817_889# a_829_889# 0.41fF
C286 a_1443_510# gnd 0.33fF
C287 a_1347_614# a_1310_617# 0.12fF
C288 a_699_455# a_711_164# 0.41fF
C289 a3_in w_310_88# 0.08fF
C290 gnd a_1472_n267# 0.21fF
C291 a_43_n236# a_36_n236# 0.41fF
C292 b1 a_733_889# 0.15fF
C293 b0 a_721_551# 0.25fF
C294 b2 a_781_889# 0.10fF
C295 w_144_n163# clk 0.08fF
C296 vdd w_405_n161# 0.17fF
C297 a_769_551# a_781_551# 0.21fF
C298 vdd w_1513_608# 0.09fF
C299 a_323_n239# a_367_n236# 0.13fF
C300 a_n85_15# vdd 0.85fF
C301 w_406_90# a_414_15# 0.10fF
C302 cin a_817_889# 0.09fF
C303 vdd a_324_12# 0.03fF
C304 a_1509_n375# a_1472_n267# 0.09fF
C305 a0 a_733_551# 0.21fF
C306 a_733_551# a3 1.49fF
C307 vdd w_1292_360# 0.08fF
C308 gnd a_n8_n239# 0.44fF
C309 a_n132_n236# a_n86_n236# 0.54fF
C310 c2 s2_out 0.09fF
C311 b0 a_n86_n236# 0.05fF
C312 a_1342_326# a_1349_326# 0.82fF
C313 a_323_n155# a_323_n239# 0.82fF
C314 w_1508_320# a_1545_326# 0.02fF
C315 cout w_985_824# 0.06fF
C316 a_1538_509# s3_out 0.41fF
C317 a_823_n105# a_712_n101# 0.06fF
C318 vdd w_29_90# 0.17fF
C319 w_812_31# a_760_37# 0.06fF
C320 a2 w_273_91# 0.06fF
C321 a_1340_37# a_1264_n67# 0.09fF
C322 vdd a_1271_510# 0.41fF
C323 vdd a_n132_n236# 0.85fF
C324 c3 w_1469_648# 0.08fF
C325 s2_out a_1521_326# 0.82fF
C326 b3 w_1341_608# 0.07fF
C327 b1 w_687_31# 0.13fF
C328 b0 vdd 1.45fF
C329 a0 w_1331_n276# 0.07fF
C330 a_771_164# a_807_164# 0.50fF
C331 w_n22_n163# a_n8_n155# 0.02fF
C332 a_759_455# w_686_449# 0.02fF
C333 a_723_455# w_883_449# 0.06fF
C334 a_711_164# w_919_379# 0.08fF
C335 clk a_n8_n239# 0.52fF
C336 a_709_889# a_721_551# 0.41fF
C337 b1 w_692_883# 0.13fF
C338 a_368_15# a_375_15# 0.41fF
C339 a_1340_37# a_1359_n68# 0.41fF
C340 vdd a_367_n236# 0.86fF
C341 a_721_551# a_733_551# 1.23fF
C342 vdd w_28_n161# 0.17fF
C343 a_1519_509# a_1482_617# 0.09fF
C344 a_1337_n375# a_1300_n267# 0.09fF
C345 a_1368_n270# vdd 0.88fF
C346 gnd a_420_n236# 0.41fF
C347 w_677_n314# n010 0.34fF
C348 a_733_551# a_745_551# 0.21fF
C349 a_711_164# b1 0.36fF
C350 a_723_455# a1 0.15fF
C351 gnd a_1477_329# 0.21fF
C352 a_712_n101# a_760_n101# 0.03fF
C353 vdd a_323_n155# 0.89fF
C354 c1 a_1512_n68# 0.09fF
C355 w_1331_n276# a_1261_n374# 0.07fF
C356 b1 c2 0.14fF
C357 a2 a_1342_326# 0.09fF
C358 a_771_455# cin 0.01fF
C359 gnd a_1303_40# 0.21fF
C360 vdd a_709_889# 0.41fF
C361 a_324_96# a_324_12# 0.82fF
C362 a_1347_614# w_1341_608# 0.21fF
C363 b0 a_724_37# 0.08fF
C364 a0 a_712_n101# 0.20fF
C365 a_1472_n267# a_1337_n270# 0.40fF
C366 s3_out gnd 0.15fF
C367 b2 c1 0.15fF
C368 a1 a_1303_40# 0.13fF
C369 b0 a_771_164# 0.01fF
C370 a_781_551# a_853_551# 0.14fF
C371 a_1342_221# a_1266_222# 0.43fF
C372 a_151_67# gnd 0.02fF
C373 a0 a_817_551# 0.23fF
C374 vdd w_n93_90# 0.17fF
C375 b3 a_1347_509# 0.09fF
C376 a_203_15# w_195_90# 0.10fF
C377 a_817_889# w_692_883# 0.11fF
C378 a_724_n101# a_736_n101# 0.26fF
C379 gnd a_414_15# 0.10fF
C380 gnd a_1340_n68# 0.52fF
C381 w_n190_n163# clk 0.08fF
C382 b2 w_686_449# 0.13fF
C383 a_1540_n270# vdd 0.88fF
C384 a1 a_1340_n68# 0.09fF
C385 w_1334_31# a_1347_37# 0.02fF
C386 gnd a_760_n101# 1.00fF
C387 a_n86_n236# a_n79_n236# 0.41fF
C388 a_1519_509# a_1347_614# 0.09fF
C389 vdd w_406_90# 0.17fF
C390 b0 a_724_n101# 0.08fF
C391 vdd w_1469_648# 0.08fF
C392 vdd w_1331_n276# 0.09fF
C393 gnd c3 0.42fF
C394 a_1310_617# a_1271_510# 0.08fF
C395 w_359_n161# a_367_n236# 0.10fF
C396 a0 w_n61_91# 0.06fF
C397 s0_out w_1503_n276# 0.21fF
C398 a1 c3 0.14fF
C399 cin w_677_n314# 0.10fF
C400 a0 gnd 1.00fF
C401 b3 a2 0.74fF
C402 b0 a_781_551# 0.09fF
C403 a3 gnd 0.54fF
C404 w_1425_253# a_1342_326# 0.24fF
C405 a_n85_15# a_n131_15# 0.54fF
C406 vdd a_1433_n374# 0.41fF
C407 w_309_n163# a_323_n239# 0.11fF
C408 a_414_15# clk 0.13fF
C409 b1 b0 8.79fF
C410 a1 a0 9.61fF
C411 a2 cin 0.73fF
C412 a1 a3 1.14fF
C413 gnd a_1361_221# 0.41fF
C414 a2 a_1305_329# 0.13fF
C415 a_1347_614# a_1347_509# 1.02fF
C416 b0 a_1300_n267# 0.13fF
C417 w_n21_88# a1_in 0.08fF
C418 a_807_455# vdd 0.41fF
C419 vdd a_1436_n67# 0.41fF
C420 vdd w_1506_31# 0.09fF
C421 gnd a_323_n239# 0.44fF
C422 gnd a_1261_n374# 0.33fF
C423 vdd a_1373_326# 0.88fF
C424 w_687_31# a_700_37# 0.02fF
C425 w_1336_320# a_1349_326# 0.02fF
C426 a_721_551# gnd 0.04fF
C427 a_n132_n236# a_n176_n239# 0.13fF
C428 a1 a_721_551# 0.35fF
C429 a2 a_733_889# 0.15fF
C430 w_902_883# a_853_889# 0.06fF
C431 vdd w_309_n163# 0.20fF
C432 a_745_551# gnd 0.21fF
C433 w_n94_n161# a_n132_n236# 0.07fF
C434 b2 w_1253_253# 0.24fF
C435 a_733_551# a_781_551# 0.77fF
C436 clk a_37_15# 0.85fF
C437 s0_out cin 0.09fF
C438 b0 a_817_889# 0.18fF
C439 a_n175_96# vdd 0.88fF
C440 a0 a_781_889# 0.21fF
C441 b1 a_733_551# 0.21fF
C442 gnd a_n86_n236# 0.10fF
C443 clk a_323_n239# 0.52fF
C444 w_1423_n36# a_1340_37# 0.24fF
C445 a_1477_329# a_1438_222# 0.08fF
C446 w_687_31# a_736_37# 0.02fF
C447 vdd w_n61_91# 0.06fF
C448 vdd a_760_37# 1.02fF
C449 w_1334_31# a_1303_40# 0.07fF
C450 a_1271_510# w_1341_608# 0.07fF
C451 a0 a_1337_n270# 0.09fF
C452 a_712_n101# a_724_37# 1.00fF
C453 vdd w_241_90# 0.17fF
C454 w_1420_n343# a_1433_n374# 0.06fF
C455 a1 vdd 1.57fF
C456 a_759_164# a_771_164# 0.21fF
C457 w_n93_90# a_n131_15# 0.07fF
C458 a_36_n236# a_n8_n239# 0.13fF
C459 w_n62_n160# a_n86_n236# 0.08fF
C460 a2 w_1336_320# 0.07fF
C461 a_723_455# w_686_449# 0.06fF
C462 a_1344_n270# vdd 0.88fF
C463 clk a_n86_n236# 0.13fF
C464 a2 w_692_883# 0.13fF
C465 w_106_n160# a_82_n236# 0.08fF
C466 w_868_14# c2 0.06fF
C467 a_817_551# a_829_551# 0.21fF
C468 w_1331_n276# a_1300_n267# 0.07fF
C469 vdd a_202_n236# 0.86fF
C470 a_1347_614# a_1354_614# 0.82fF
C471 vdd w_n62_n160# 0.06fF
C472 a_414_15# a_421_15# 0.41fF
C473 s3_out a_1550_614# 0.82fF
C474 vdd clk 1.34fF
C475 b2_in a_158_n239# 0.07fF
C476 a_712_n101# a_724_n101# 0.58fF
C477 a_1261_n374# a_1337_n270# 0.09fF
C478 gnd a_1266_222# 0.33fF
C479 a_711_164# a2 0.26fF
C480 gnd a_210_15# 0.41fF
C481 a_203_15# a_159_12# 0.13fF
C482 a2 c2 0.14fF
C483 a_771_455# b0 0.01fF
C484 gnd s2_out 0.15fF
C485 a_255_n236# a_248_n236# 0.41fF
C486 a_724_37# a_760_37# 0.82fF
C487 vdd s1_out 0.05fF
C488 cin n010 0.00fF
C489 a_n175_96# a_n175_12# 0.82fF
C490 a_368_15# a_324_12# 0.13fF
C491 cin w_1503_n276# 0.07fF
C492 b1 a_712_n101# 0.14fF
C493 a1 a_724_37# 0.01fF
C494 a_829_551# gnd 0.21fF
C495 a_1516_n270# vdd 0.88fF
C496 a1 a_771_164# 0.01fF
C497 a0 a_723_164# 0.15fF
C498 c3 c1 0.10fF
C499 a_781_551# a_817_551# 0.83fF
C500 vdd a_1378_614# 0.88fF
C501 gnd a_n124_15# 0.41fF
C502 a_1305_329# a_1342_326# 0.12fF
C503 vdd w_n189_88# 0.20fF
C504 a_1347_509# a_1271_510# 0.43fF
C505 a0 c1 0.15fF
C506 a3 c1 0.15fF
C507 a_151_67# w_145_88# 0.08fF
C508 a_1514_221# a_1342_326# 0.09fF
C509 a_n175_12# gnd 0.44fF
C510 a_769_889# w_692_883# 0.02fF
C511 w_145_88# a_159_96# 0.02fF
C512 a_83_15# w_75_90# 0.10fF
C513 gnd a_724_n101# 0.05fF
C514 a2 w_1292_360# 0.08fF
C515 b0 w_844_449# 0.06fF
C516 a0 w_686_449# 0.13fF
C517 vdd a_1337_n270# 0.14fF
C518 vdd w_310_88# 0.20fF
C519 a1 a_724_n101# 0.01fF
C520 w_1506_31# a_1519_37# 0.02fF
C521 vdd w_1297_648# 0.08fF
C522 w_309_n163# b3_in 0.08fF
C523 gnd a_1310_617# 0.21fF
C524 gnd b0_in 0.02fF
C525 a_690_n370# n010 0.25fF
C526 w_359_n161# clk 0.07fF
C527 b0 w_677_n314# 0.10fF
C528 b1 gnd 0.94fF
C529 a0 a_853_889# 0.09fF
C530 b2 c3 0.14fF
C531 a1 a_781_551# 0.09fF
C532 w_1508_320# a_1342_326# 0.07fF
C533 a_n175_12# clk 0.52fF
C534 b2 a0 1.10fF
C535 b3 cin 2.20fF
C536 a1 b1 6.23fF
C537 a2 b0 2.20fF
C538 b2 a3 0.86fF
C539 a_83_15# a_37_15# 0.54fF
C540 gnd a_1300_n267# 0.21fF
C541 gnd b3_in 0.02fF
C542 a_1443_510# s3_out 0.09fF
C543 w_n21_88# clk 0.08fF
C544 a2 a_1342_221# 0.09fF
C545 a_759_455# vdd 0.41fF
C546 a_1337_n375# a_1356_n375# 0.08fF
C547 w_1430_541# a_1347_614# 0.24fF
C548 vdd w_1334_31# 0.09fF
C549 vdd a_690_n308# 0.41fF
C550 gnd a_89_n236# 0.41fF
C551 vdd a_1438_222# 0.41fF
C552 w_812_31# a_823_n105# 0.07fF
C553 a_n175_12# w_n189_88# 0.11fF
C554 w_1336_320# a_1342_326# 0.21fF
C555 b3 a_413_n236# 0.05fF
C556 w_74_n161# a_36_n236# 0.07fF
C557 gnd a_n176_n239# 0.44fF
C558 a_1519_509# a_1538_509# 0.08fF
C559 vdd c1 1.48fF
C560 b2 a_721_551# 0.41fF
C561 a_1443_510# c3 0.56fF
C562 w_n22_n163# clk 0.08fF
C563 b3 a_1347_614# 0.09fF
C564 a_1347_614# a_1482_617# 0.40fF
C565 a_709_551# gnd 0.21fF
C566 vdd w_240_n161# 0.17fF
C567 vdd a_1550_614# 0.88fF
C568 vdd w_n140_n161# 0.17fF
C569 clk a_n131_15# 0.86fF
C570 a_368_15# w_406_90# 0.07fF
C571 w_310_88# a_324_96# 0.02fF
C572 a1 a_817_889# 0.09fF
C573 b1 a_781_889# 0.10fF
C574 cin a_733_889# 0.08fF
C575 vdd a_249_15# 0.86fF
C576 a2 a_733_551# 0.21fF
C577 a_771_455# a_807_455# 1.04fF
C578 vdd w_686_449# 0.17fF
C579 a_1340_37# a_1436_n67# 0.20fF
C580 a_83_15# vdd 0.86fF
C581 a_711_164# a_699_164# 0.21fF
C582 w_1420_n343# a_1337_n270# 0.24fF
C583 gnd a_248_n236# 0.10fF
C584 w_1506_31# a_1340_37# 0.07fF
C585 c2 a_1342_326# 0.57fF
C586 clk a_n176_n239# 0.52fF
C587 s0_out a_1528_n375# 0.41fF
C588 vdd a_853_889# 0.41fF
C589 a_1438_222# s2_out 0.09fF
C590 a_1310_617# w_1297_648# 0.06fF
C591 a_700_37# a_712_n101# 0.41fF
C592 vdd w_145_88# 0.20fF
C593 a_1436_n67# a_1475_40# 0.08fF
C594 w_1506_31# a_1475_40# 0.07fF
C595 b2 vdd 1.38fF
C596 s1_out a_1519_37# 0.82fF
C597 w_n139_90# clk 0.07fF
C598 a_829_889# w_692_883# 0.02fF
C599 a3 w_941_883# 0.06fF
C600 a_723_164# a_771_164# 0.50fF
C601 a_699_455# w_686_449# 0.02fF
C602 a_248_n236# a_202_n236# 0.54fF
C603 cin w_687_31# 0.06fF
C604 b3 w_692_883# 0.14fF
C605 a_1300_n267# a_1337_n270# 0.12fF
C606 clk a_248_n236# 0.13fF
C607 a_807_455# w_844_449# 0.06fF
C608 cin w_692_883# 0.06fF
C609 vdd a_36_n236# 0.86fF
C610 a_1519_509# gnd 0.52fF
C611 w_1336_320# a_1305_329# 0.07fF
C612 w_360_90# clk 0.07fF
C613 a_781_889# a_817_889# 1.20fF
C614 w_868_14# a_712_n101# 0.08fF
C615 cin w_1459_n236# 0.08fF
C616 vdd w_144_n163# 0.20fF
C617 gnd a_1340_37# 0.26fF
C618 w_1513_608# a_1526_614# 0.02fF
C619 a_1303_40# a_1340_n68# 0.09fF
C620 b2 a_1266_222# 0.20fF
C621 b3 c2 0.14fF
C622 a_771_455# a1 0.01fF
C623 a_711_164# cin 0.19fF
C624 a_723_455# a0 0.15fF
C625 s0_out a_1540_n270# 0.82fF
C626 a1 a_1340_37# 0.09fF
C627 w_144_n163# a_158_n155# 0.02fF
C628 b1 w_1334_31# 0.07fF
C629 vdd a_1347_37# 0.88fF
C630 b0 n010 0.01fF
C631 gnd a_735_164# 0.21fF
C632 a_721_551# w_941_883# 0.06fF
C633 a_714_n308# w_749_n314# 0.06fF
C634 gnd a_1475_40# 0.21fF
C635 b1 a_723_164# 0.15fF
C636 vdd a_745_889# 0.41fF
C637 vdd a_1443_510# 0.41fF
C638 a_1378_614# w_1341_608# 0.02fF
C639 s3_out c3 0.09fF
C640 a_1347_509# gnd 0.52fF
C641 vdd w_1253_253# 0.06fF
C642 vdd a_1472_n267# 0.44fF
C643 b1 c1 0.15fF
C644 cin a_807_164# 0.09fF
C645 a_733_889# w_692_883# 0.07fF
C646 a_1342_221# a_1342_326# 1.02fF
C647 a_1514_221# c2 0.09fF
C648 s0_out a_1433_n374# 0.09fF
C649 gnd a_44_15# 0.41fF
C650 w_1513_608# a_1482_617# 0.07fF
C651 a_1533_221# s2_out 0.41fF
C652 vdd a_n8_n239# 0.03fF
C653 b0 w_1287_n236# 0.08fF
C654 gnd a_1531_n68# 0.41fF
C655 b1 w_686_449# 0.13fF
C656 a2 w_883_449# 0.06fF
C657 w_1258_541# a3 0.24fF
C658 s1_out a_1340_37# 0.09fF
C659 a3 a_414_15# 0.05fF
C660 cout gnd 0.21fF
C661 b3 a_1271_510# 0.56fF
C662 a2 gnd 0.78fF
C663 b2 a_781_551# 0.09fF
C664 w_1292_360# a_1305_329# 0.06fF
C665 w_1253_253# a_1266_222# 0.06fF
C666 w_1464_360# a_1477_329# 0.06fF
C667 w_1508_320# c2 0.07fF
C668 a_368_15# clk 0.85fF
C669 a2 a1 6.02fF
C670 b3 b0 0.91fF
C671 b2 b1 7.89fF
C672 s1_out a_1475_40# 0.12fF
C673 a0 c3 0.14fF
C674 a3 c3 0.14fF
C675 w_1508_320# a_1521_326# 0.02fF
C676 a_n7_12# a1_in 0.07fF
C677 w_405_n161# a_413_n236# 0.10fF
C678 b0 cin 1.67fF
C679 gnd b2_in 0.02fF
C680 a0 a3 1.14fF
C681 gnd a0_in 0.02fF
C682 a_1540_n270# w_1503_n276# 0.02fF
C683 w_1513_608# a_1347_614# 0.07fF
C684 w_195_90# clk 0.07fF
C685 w_75_90# a_37_15# 0.07fF
C686 s1_out a_1531_n68# 0.41fF
C687 vdd a_1477_329# 0.44fF
C688 vdd w_n190_n163# 0.20fF
C689 w_240_n161# a_248_n236# 0.10fF
C690 a_1342_221# a_1305_329# 0.09fF
C691 w_812_31# a_724_37# 0.06fF
C692 vdd a_1303_40# 0.44fF
C693 a0 a_1261_n374# 0.20fF
C694 s0_out gnd 0.13fF
C695 w_782_n313# c1 0.06fF
C696 w_1503_n276# a_1433_n374# 0.07fF
C697 a_817_889# a_853_889# 1.79fF
C698 w_194_n161# a_202_n236# 0.10fF
C699 a_1347_614# a_1271_510# 0.09fF
C700 vdd s3_out 0.05fF
C701 a2 a_781_889# 0.10fF
C702 a0 a_721_551# 0.25fF
C703 b0 a_733_889# 0.15fF
C704 vdd a_159_96# 0.89fF
C705 w_194_n161# clk 0.07fF
C706 a_721_551# a3 0.24fF
C707 vdd w_437_n160# 0.06fF
C708 s0_out a_1509_n375# 1.02fF
C709 vdd w_1258_541# 0.06fF
C710 a_759_455# a_771_455# 0.41fF
C711 a_413_n236# a_367_n236# 0.54fF
C712 a_n7_96# vdd 0.89fF
C713 w_438_91# a_414_15# 0.08fF
C714 w_1334_31# a_1340_37# 0.21fF
C715 vdd a_414_15# 0.86fF
C716 cin a_733_551# 0.10fF
C717 gnd a_82_n236# 0.10fF
C718 b2 a_248_n236# 0.05fF
C719 a_1477_329# s2_out 0.12fF
C720 a_1342_326# a_1373_326# 0.82fF
C721 a_1366_509# a_1347_509# 0.08fF
C722 a_823_n105# a_724_37# 0.01fF
C723 vdd w_75_90# 0.17fF
C724 vdd c3 1.01fF
C725 a_1340_37# c1 0.57fF
C726 w_1462_71# c1 0.08fF
C727 a_1482_617# w_1469_648# 0.06fF
C728 a_723_164# a_735_164# 0.21fF
C729 w_n189_88# a0_in 0.08fF
C730 a1 w_1290_71# 0.08fF
C731 b0 w_687_31# 0.06fF
C732 a0 vdd 2.64fF
C733 w_438_91# a3 0.06fF
C734 vdd a3 1.33fF
C735 w_n22_n163# a_n8_n239# 0.11fF
C736 a_771_455# w_686_449# 0.06fF
C737 a_1337_n375# b0 0.09fF
C738 clk a_82_n236# 0.13fF
C739 b0 w_692_883# 0.06fF
C740 c1 a_1475_40# 0.13fF
C741 s0_out a_1516_n270# 0.82fF
C742 a_1340_37# a_1512_n68# 0.09fF
C743 cin a_1433_n374# 0.56fF
C744 a_769_889# a_781_889# 0.41fF
C745 a_1356_n375# gnd 0.41fF
C746 vdd w_74_n161# 0.17fF
C747 a_823_n105# a_724_n101# 0.08fF
C748 gnd n010 0.26fF
C749 w_677_n314# a_690_n308# 0.02fF
C750 vdd a_37_15# 0.86fF
C751 w_902_883# a_817_889# 0.06fF
C752 a_723_455# b1 0.15fF
C753 a_711_164# b0 0.26fF
C754 gnd a_1342_326# 0.26fF
C755 gnd a_375_15# 0.41fF
C756 vdd a_323_n239# 0.03fF
C757 w_n190_n163# b0_in 0.08fF
C758 vdd a_1261_n374# 0.41fF
C759 a_1475_40# a_1512_n68# 0.09fF
C760 gnd a_699_164# 0.21fF
C761 a_n85_15# a_n78_15# 0.41fF
C762 b0 c2 0.14fF
C763 a_807_455# cin 0.06fF
C764 s0_out a_1337_n270# 0.09fF
C765 gnd a_1264_n67# 0.33fF
C766 a0 a_724_37# 0.15fF
C767 cin a_712_n101# 0.14fF
C768 vdd w_1464_360# 0.08fF
C769 w_1506_31# a_1543_37# 0.02fF
C770 a_374_n236# a_367_n236# 0.41fF
C771 b1 a_1303_40# 0.40fF
C772 a2 c1 0.15fF
C773 a0 a_771_164# 0.01fF
C774 a1 a_1264_n67# 0.56fF
C775 a_709_889# w_692_883# 0.02fF
C776 a_1512_n68# a_1531_n68# 0.08fF
C777 b2 w_272_n160# 0.06fF
C778 gnd a_159_12# 0.44fF
C779 cin a_817_551# 0.12fF
C780 a_203_15# w_241_90# 0.07fF
C781 a_n7_96# w_n21_88# 0.02fF
C782 a_724_n101# a_760_n101# 0.56fF
C783 a_n7_12# gnd 0.44fF
C784 vdd a_n86_n236# 0.85fF
C785 a2 a_249_15# 0.05fF
C786 gnd a_1359_n68# 0.41fF
C787 a2 w_686_449# 0.06fF
C788 w_919_379# c3 0.06fF
C789 b1 a_1340_n68# 0.09fF
C790 a_1347_37# a_1340_37# 0.82fF
C791 gnd a_209_n236# 0.41fF
C792 w_1334_31# a_1371_37# 0.02fF
C793 a_1519_509# a_1443_510# 0.43fF
C794 vdd w_438_91# 0.06fF
C795 a0 a_724_n101# 0.15fF
C796 b3 gnd 0.63fF
C797 w_405_n161# a_367_n236# 0.07fF
C798 gnd a_1482_617# 0.21fF
C799 w_n190_n163# a_n176_n239# 0.11fF
C800 a_1516_n270# w_1503_n276# 0.02fF
C801 a_203_15# clk 0.85fF
C802 a1 w_107_91# 0.06fF
C803 a_159_12# clk 0.52fF
C804 b1 c3 0.14fF
C805 b3 a1 0.99fF
C806 b2 a2 4.39fF
C807 vdd a_158_n155# 0.89fF
C808 cin gnd 0.26fF
C809 a0 a_781_551# 0.18fF
C810 a3 a_1310_617# 0.40fF
C811 w_1425_253# a_1438_222# 0.06fF
C812 a_n7_12# clk 0.52fF
C813 b1 a0 1.52fF
C814 a1 cin 1.10fF
C815 a_202_n236# a_209_n236# 0.41fF
C816 gnd b1_in 0.02fF
C817 b1 a3 0.85fF
C818 a_1356_n375# a_1337_n270# 0.41fF
C819 cin a_1509_n375# 0.09fF
C820 gnd a_1305_329# 0.21fF
C821 gnd a_1514_221# 0.52fF
C822 a_699_455# vdd 0.41fF
C823 a0 a_1300_n267# 0.40fF
C824 w_749_n314# n010 0.06fF
C825 w_1503_n276# a_1337_n270# 0.07fF
C826 vdd a_1266_222# 0.41fF
C827 vdd w_1251_n36# 0.06fF
C828 gnd a_413_n236# 0.10fF
C829 vdd s2_out 0.05fF
C830 w_687_31# a_712_n101# 0.09fF
C831 a_n85_15# w_n93_90# 0.10fF
C832 w_1336_320# a_1373_326# 0.02fF
C833 a_690_n370# gnd 0.21fF
C834 a_1347_614# gnd 0.26fF
C835 w_144_n163# b2_in 0.08fF
C836 a_714_n308# a0 0.08fF
C837 b1 a_721_551# 0.25fF
C838 a1 a_733_889# 0.15fF
C839 w_273_91# a_249_15# 0.08fF
C840 vdd w_359_n161# 0.17fF
C841 a_769_551# gnd 0.21fF
C842 a_723_455# a_771_455# 0.97fF
C843 a_1300_n267# a_1261_n374# 0.08fF
C844 s1_out a_1543_37# 0.82fF
C845 a_323_n239# b3_in 0.07fF
C846 a0 a_817_889# 0.18fF
C847 a_n175_12# vdd 0.03fF
C848 cin a_781_889# 0.10fF
C849 vdd a_324_96# 0.89fF
C850 b0 a_733_551# 0.21fF
C851 n010 a_690_n308# 0.41fF
C852 vdd w_919_379# 0.06fF
C853 clk a_413_n236# 0.13fF
C854 w_1423_n36# a_1436_n67# 0.06fF
C855 vdd w_1420_n343# 0.06fF
C856 a_1342_326# a_1438_222# 0.20fF
C857 a_712_n101# c2 0.05fF
C858 a_1519_509# s3_out 1.02fF
C859 w_687_31# a_760_37# 0.03fF
C860 vdd w_n21_88# 0.20fF
C861 a_1340_37# a_1303_40# 0.12fF
C862 w_1334_31# a_1264_n67# 0.07fF
C863 b3 w_1297_648# 0.08fF
C864 vdd a_1310_617# 0.44fF
C865 n010 c1 0.05fF
C866 cin a_1337_n270# 0.57fF
C867 a1 w_687_31# 0.13fF
C868 a_1337_n375# gnd 0.52fF
C869 b1 vdd 1.34fF
C870 a3 w_1341_608# 0.07fF
C871 gnd a_158_n239# 0.44fF
C872 a_36_n236# a_82_n236# 0.54fF
C873 b0 w_1331_n276# 0.07fF
C874 a_711_164# w_883_449# 0.06fF
C875 a_735_455# w_686_449# 0.02fF
C876 a1 w_692_883# 0.13fF
C877 a_1340_37# a_1340_n68# 1.02fF
C878 a_817_551# a_853_551# 0.78fF
C879 vdd a_1300_n267# 0.44fF
C880 vdd a_1545_326# 0.88fF
C881 a_733_889# a_781_889# 1.27fF
C882 a_721_551# a_709_551# 0.21fF
C883 a_1347_614# a_1378_614# 0.82fF
C884 vdd w_n22_n163# 0.20fF
C885 a_1519_509# c3 0.09fF
C886 s0_out a_1472_n267# 0.12fF
C887 a_711_164# gnd 0.04fF
C888 vdd a_n131_15# 0.85fF
C889 gnd a_374_n236# 0.41fF
C890 a_1368_n270# w_1331_n276# 0.02fF
C891 a_202_n236# a_158_n239# 0.13fF
C892 a_711_164# a1 0.28fF
C893 gnd c2 0.42fF
C894 gnd a_256_15# 0.41fF
C895 a_203_15# a_249_15# 0.54fF
C896 clk a_158_n239# 0.52fF
C897 b2 a_1342_326# 0.09fF
C898 a1 c2 0.14fF
C899 a_771_455# a0 0.01fF
C900 w_n94_n161# a_n86_n236# 0.10fF
C901 vdd a_1519_37# 0.88fF
C902 b1 w_1251_n36# 0.24fF
C903 a_714_n308# vdd 0.41fF
C904 gnd a_807_164# 0.23fF
C905 a_368_15# a_414_15# 0.54fF
C906 vdd a_n176_n239# 0.03fF
C907 b0 a_712_n101# 0.14fF
C908 a_853_551# gnd 0.21fF
C909 b1 a_771_164# 0.01fF
C910 b3 c1 0.15fF
C911 cin a_723_164# 0.08fF
C912 vdd w_n94_n161# 0.17fF
C913 b0 a_817_551# 0.23fF
C914 gnd a_n78_15# 0.41fF
C915 vdd w_n139_90# 0.17fF
C916 a1 a_853_551# 0.09fF
C917 cin c1 0.16fF
C918 a_n85_15# w_n61_91# 0.08fF
C919 w_145_88# a_159_12# 0.11fF
C920 a_n85_15# gnd 0.10fF
C921 a_1545_326# s2_out 0.82fF
C922 a_781_889# w_692_883# 0.19fF
C923 a_1514_221# a_1438_222# 0.43fF
C924 gnd a_324_12# 0.44fF
C925 a0 w_1248_n343# 0.24fF
C926 a_1347_509# a3 0.09fF
C927 w_n190_n163# a_n176_n155# 0.02fF
C928 vdd a_248_n236# 0.86fF
C929 a_83_15# w_107_91# 0.08fF
C930 gnd a_736_n101# 0.21fF
C931 a_1366_509# a_1347_614# 0.41fF
C932 cin w_686_449# 0.06fF
C933 vdd w_360_90# 0.17fF
C934 vdd w_1341_608# 0.09fF
C935 vdd w_782_n313# 0.10fF
C936 a_714_n370# n010 0.64fF
C937 gnd a_1271_510# 0.33fF
C938 a_1337_n375# a_1337_n270# 1.02fF
C939 a_n124_15# a_n131_15# 0.41fF
C940 b3 b2 5.56fF
C941 a0 w_677_n314# 0.21fF
C942 b0 gnd 1.42fF
C943 a2 c3 0.14fF
C944 b1 a_781_551# 0.09fF
C945 w_1508_320# a_1438_222# 0.07fF
C946 w_309_n163# a_323_n155# 0.02fF
C947 a_n175_12# a_n131_15# 0.13fF
C948 a_n85_15# clk 0.13fF
C949 a_44_15# a_37_15# 0.41fF
C950 w_1503_n276# a_1472_n267# 0.07fF
C951 a_324_12# clk 0.52fF
C952 w_1248_n343# a_1261_n374# 0.06fF
C953 b2 cin 0.61fF
C954 a1 b0 2.49fF
C955 a2 a0 1.34fF
C956 a2 a3 3.43fF
C957 a_1528_n375# Gnd 0.02fF
C958 a_1509_n375# Gnd 0.26fF
C959 a_1356_n375# Gnd 0.02fF
C960 a_1337_n375# Gnd 0.26fF
C961 a_1540_n270# Gnd 0.00fF
C962 a_1516_n270# Gnd 0.00fF
C963 s0_out Gnd 0.64fF
C964 a_714_n370# Gnd 0.24fF
C965 a_690_n370# Gnd 0.04fF
C966 a_1368_n270# Gnd 0.00fF
C967 a_1344_n270# Gnd 0.00fF
C968 a_714_n308# Gnd 0.15fF
C969 a_690_n308# Gnd 0.00fF
C970 n010 Gnd 3.19fF
C971 a_420_n236# Gnd 0.02fF
C972 a_374_n236# Gnd 0.02fF
C973 a_1433_n374# Gnd 1.23fF
C974 a_1337_n270# Gnd 2.69fF
C975 a_1472_n267# Gnd 0.76fF
C976 a_1261_n374# Gnd 1.23fF
C977 a_1300_n267# Gnd 0.76fF
C978 a_255_n236# Gnd 0.02fF
C979 a_209_n236# Gnd 0.02fF
C980 a_760_n101# Gnd 0.24fF
C981 a_736_n101# Gnd 0.02fF
C982 a_724_n101# Gnd 0.65fF
C983 a_700_n101# Gnd 0.02fF
C984 a_1531_n68# Gnd 0.02fF
C985 a_1512_n68# Gnd 0.26fF
C986 a_1359_n68# Gnd 0.02fF
C987 a_1340_n68# Gnd 0.26fF
C988 a_1543_37# Gnd 0.00fF
C989 a_1519_37# Gnd 0.00fF
C990 s1_out Gnd 0.64fF
C991 a_1371_37# Gnd 0.00fF
C992 a_1347_37# Gnd 0.00fF
C993 a_413_n236# Gnd 0.75fF
C994 a_323_n239# Gnd 0.25fF
C995 a_323_n155# Gnd 0.00fF
C996 a_89_n236# Gnd 0.02fF
C997 a_43_n236# Gnd 0.02fF
C998 a_248_n236# Gnd 0.75fF
C999 a_158_n155# Gnd 0.00fF
C1000 a_n79_n236# Gnd 0.02fF
C1001 a_n125_n236# Gnd 0.02fF
C1002 a_82_n236# Gnd 0.75fF
C1003 a_n8_n239# Gnd 0.18fF
C1004 a_n8_n155# Gnd 0.00fF
C1005 a_n86_n236# Gnd 0.75fF
C1006 a_n176_n239# Gnd 0.18fF
C1007 a_n176_n155# Gnd 0.00fF
C1008 a_367_n236# Gnd 1.01fF
C1009 b3_in Gnd 0.34fF
C1010 a_202_n236# Gnd 1.01fF
C1011 b2_in Gnd 0.34fF
C1012 a_36_n236# Gnd 1.01fF
C1013 b1_in Gnd 0.28fF
C1014 a_n132_n236# Gnd 1.01fF
C1015 b0_in Gnd 0.28fF
C1016 a_760_37# Gnd 0.26fF
C1017 a_736_37# Gnd 0.00fF
C1018 a_724_37# Gnd 0.73fF
C1019 a_712_n101# Gnd 1.83fF
C1020 a_700_37# Gnd 0.00fF
C1021 a_421_15# Gnd 0.02fF
C1022 a_375_15# Gnd 0.02fF
C1023 a_823_n105# Gnd 0.69fF
C1024 a_256_15# Gnd 0.02fF
C1025 a_210_15# Gnd 0.02fF
C1026 a_1436_n67# Gnd 1.23fF
C1027 a_1340_37# Gnd 2.69fF
C1028 a_1475_40# Gnd 0.76fF
C1029 c1 Gnd 19.81fF
C1030 a_1264_n67# Gnd 1.23fF
C1031 a_1303_40# Gnd 0.76fF
C1032 a_807_164# Gnd 0.22fF
C1033 a_771_164# Gnd 1.17fF
C1034 a_759_164# Gnd 0.02fF
C1035 a_735_164# Gnd 0.02fF
C1036 a_723_164# Gnd 1.01fF
C1037 a_699_164# Gnd 0.02fF
C1038 a_414_15# Gnd 0.75fF
C1039 a_324_12# Gnd 0.48fF
C1040 a_324_96# Gnd 0.00fF
C1041 a_90_15# Gnd 0.02fF
C1042 a_44_15# Gnd 0.02fF
C1043 a_249_15# Gnd 0.75fF
C1044 a_159_12# Gnd 0.48fF
C1045 a_159_96# Gnd 0.00fF
C1046 a_n78_15# Gnd 0.02fF
C1047 a_n124_15# Gnd 0.02fF
C1048 a_83_15# Gnd 0.75fF
C1049 a_n7_12# Gnd 0.48fF
C1050 a_n7_96# Gnd 0.00fF
C1051 a_n85_15# Gnd 0.75fF
C1052 a_n175_12# Gnd 0.48fF
C1053 a_n175_96# Gnd 0.00fF
C1054 a_368_15# Gnd 1.01fF
C1055 a3_in Gnd 0.21fF
C1056 a_203_15# Gnd 1.01fF
C1057 a_151_67# Gnd 0.06fF
C1058 a_37_15# Gnd 1.01fF
C1059 a1_in Gnd 0.15fF
C1060 a_n131_15# Gnd 1.01fF
C1061 clk Gnd 0.09fF
C1062 a0_in Gnd 0.34fF
C1063 a_1533_221# Gnd 0.02fF
C1064 a_1514_221# Gnd 0.26fF
C1065 a_1361_221# Gnd 0.02fF
C1066 a_1342_221# Gnd 0.26fF
C1067 a_1545_326# Gnd 0.00fF
C1068 a_1521_326# Gnd 0.00fF
C1069 s2_out Gnd 0.63fF
C1070 a_1373_326# Gnd 0.00fF
C1071 a_1349_326# Gnd 0.00fF
C1072 a_1438_222# Gnd 1.23fF
C1073 a_1342_326# Gnd 2.69fF
C1074 a_1477_329# Gnd 0.76fF
C1075 c2 Gnd 14.66fF
C1076 a_1266_222# Gnd 1.23fF
C1077 a_1305_329# Gnd 0.76fF
C1078 a_807_455# Gnd 0.20fF
C1079 a_771_455# Gnd 1.16fF
C1080 a_759_455# Gnd 0.00fF
C1081 a_735_455# Gnd 0.00fF
C1082 a_723_455# Gnd 0.92fF
C1083 a_711_164# Gnd 3.38fF
C1084 a_699_455# Gnd 0.00fF
C1085 a_1538_509# Gnd 0.02fF
C1086 a_1519_509# Gnd 0.26fF
C1087 a_1366_509# Gnd 0.02fF
C1088 a_1347_509# Gnd 0.26fF
C1089 a_1550_614# Gnd 0.00fF
C1090 a_1526_614# Gnd 0.00fF
C1091 s3_out Gnd 0.63fF
C1092 a_853_551# Gnd 0.30fF
C1093 a_829_551# Gnd 0.02fF
C1094 a_817_551# Gnd 0.89fF
C1095 a_781_551# Gnd 1.29fF
C1096 a_769_551# Gnd 0.02fF
C1097 a_745_551# Gnd 0.02fF
C1098 a_733_551# Gnd 2.00fF
C1099 a_709_551# Gnd 0.02fF
C1100 a_1378_614# Gnd 0.00fF
C1101 a_1354_614# Gnd 0.00fF
C1102 a_1443_510# Gnd 1.23fF
C1103 a_1347_614# Gnd 2.69fF
C1104 a_1482_617# Gnd 0.76fF
C1105 c3 Gnd 10.13fF
C1106 a_1271_510# Gnd 1.23fF
C1107 a_1310_617# Gnd 0.76fF
C1108 gnd Gnd 0.17fF
C1109 cout Gnd 0.10fF
C1110 a_853_889# Gnd 0.23fF
C1111 a_829_889# Gnd 0.00fF
C1112 a_817_889# Gnd 0.59fF
C1113 a_781_889# Gnd 0.98fF
C1114 a_769_889# Gnd 0.00fF
C1115 a_745_889# Gnd 0.00fF
C1116 a_733_889# Gnd 1.46fF
C1117 a_721_551# Gnd 4.42fF
C1118 a_709_889# Gnd 0.00fF
C1119 vdd Gnd 30.98fF
C1120 cin Gnd 25.39fF
C1121 a0 Gnd 58.07fF
C1122 b0 Gnd 55.49fF
C1123 b1 Gnd 51.60fF
C1124 a1 Gnd 55.50fF
C1125 a2 Gnd 50.88fF
C1126 b2 Gnd 47.22fF
C1127 b3 Gnd 39.18fF
C1128 a3 Gnd 42.69fF
C1129 w_1420_n343# Gnd 1.25fF
C1130 w_1248_n343# Gnd 1.25fF
C1131 w_1503_n276# Gnd 5.54fF
C1132 w_1459_n236# Gnd 1.25fF
C1133 w_1331_n276# Gnd 5.54fF
C1134 w_782_n313# Gnd 1.25fF
C1135 w_749_n314# Gnd 1.38fF
C1136 w_677_n314# Gnd 3.51fF
C1137 w_1287_n236# Gnd 1.25fF
C1138 w_437_n160# Gnd 1.46fF
C1139 w_405_n161# Gnd 2.53fF
C1140 w_359_n161# Gnd 2.53fF
C1141 w_309_n163# Gnd 3.68fF
C1142 w_272_n160# Gnd 1.46fF
C1143 w_240_n161# Gnd 2.53fF
C1144 w_194_n161# Gnd 2.53fF
C1145 w_144_n163# Gnd 0.02fF
C1146 w_106_n160# Gnd 1.46fF
C1147 w_74_n161# Gnd 2.53fF
C1148 w_28_n161# Gnd 2.53fF
C1149 w_n22_n163# Gnd 3.68fF
C1150 w_n62_n160# Gnd 1.46fF
C1151 w_n94_n161# Gnd 2.53fF
C1152 w_n140_n161# Gnd 2.53fF
C1153 w_n190_n163# Gnd 3.68fF
C1154 w_1423_n36# Gnd 1.25fF
C1155 w_1251_n36# Gnd 1.25fF
C1156 w_1506_31# Gnd 5.54fF
C1157 w_1462_71# Gnd 1.25fF
C1158 w_1334_31# Gnd 5.54fF
C1159 w_868_14# Gnd 1.25fF
C1160 w_1290_71# Gnd 1.25fF
C1161 w_812_31# Gnd 1.25fF
C1162 w_687_31# Gnd 5.64fF
C1163 w_438_91# Gnd 1.46fF
C1164 w_406_90# Gnd 2.53fF
C1165 w_360_90# Gnd 2.53fF
C1166 w_310_88# Gnd 0.04fF
C1167 w_273_91# Gnd 1.46fF
C1168 w_241_90# Gnd 2.53fF
C1169 w_195_90# Gnd 2.53fF
C1170 w_145_88# Gnd 3.68fF
C1171 w_107_91# Gnd 1.46fF
C1172 w_75_90# Gnd 2.53fF
C1173 w_29_90# Gnd 2.53fF
C1174 w_n21_88# Gnd 3.68fF
C1175 w_n61_91# Gnd 1.46fF
C1176 w_n93_90# Gnd 2.53fF
C1177 w_n139_90# Gnd 2.53fF
C1178 w_n189_88# Gnd 3.68fF
C1179 w_1425_253# Gnd 1.25fF
C1180 w_1253_253# Gnd 1.25fF
C1181 w_1508_320# Gnd 5.54fF
C1182 w_1464_360# Gnd 1.25fF
C1183 w_1336_320# Gnd 5.54fF
C1184 w_1292_360# Gnd 1.25fF
C1185 w_919_379# Gnd 1.25fF
C1186 w_883_449# Gnd 1.33fF
C1187 w_844_449# Gnd 1.33fF
C1188 w_686_449# Gnd 7.72fF
C1189 w_1430_541# Gnd 1.25fF
C1190 w_1258_541# Gnd 1.25fF
C1191 w_1513_608# Gnd 5.54fF
C1192 w_1469_648# Gnd 1.25fF
C1193 w_1341_608# Gnd 5.54fF
C1194 w_1297_648# Gnd 1.25fF
C1195 w_985_824# Gnd 1.25fF
C1196 w_941_883# Gnd 1.33fF
C1197 w_902_883# Gnd 1.33fF
C1198 w_692_883# Gnd 10.49fF

.tran 10n 1u

.control
set hcopypscolor = 1 
set color0=white
set color1=black
run


plot V(a3) V(b3)+2 V(c3)+4 V(s3_out)+6 V(cout)+8
*plot V(a0) V(b0)+2 V(a1)+4 V(b1)+6 
*plot V(a2) V(b2)+2 V(a3)+4 V(b3)+6 V(cout)+8
*plot V(a3) V(b3)+2 V(cout)+4
.endc
.end