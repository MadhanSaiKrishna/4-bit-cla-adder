.subckt carry_one c1 A0 B0 Cin vdd gnd

.param width_P = 40*LAMBDA
.param width_N = 20*LAMBDA

* M1 n1 A0 gnd gnd CMOSN W={width_N} L={2*LAMBDA}
* +AS={5*width_N*LAMBDA} PS={10*LAMBDA+width_N}
* +AD={5*width_N*LAMBDA} PD={10*LAMBDA+width_N}

* M2 n2 B0 n1 n1 CMOSN W={width_N} L={2*LAMBDA}
* +AS={5*width_N*LAMBDA} PS={10*LAMBDA+width_N}
* +AD={5*width_N*LAMBDA} PD={10*LAMBDA+width_N}

* M3 n2 B0 n3 n3 CMOSP W={width_P} L={2*LAMBDA}
* +AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
* +AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

* M4 n3 A0 vdd vdd CMOSP W={width_P} L={2*LAMBDA}
* +AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
* +AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

* M5 n2 A0 n4 n4 CMOSN W={width_N} L={2*LAMBDA}
* +AS={5*width_N*LAMBDA} PS={10*LAMBDA+width_N}
* +AD={5*width_N*LAMBDA} PD={10*LAMBDA+width_N}

* M6 n2 B0 n4 n4 CMOSN W={width_N} L={2*LAMBDA}
* +AS={5*width_N*LAMBDA} PS={10*LAMBDA+width_N}
* +AD={5*width_N*LAMBDA} PD={10*LAMBDA+width_N}

* M7 n4 Cin gnd gnd CMOSN W={width_N} L={2*LAMBDA}
* +AS={5*width_N*LAMBDA} PS={10*LAMBDA+width_N}
* +AD={5*width_N*LAMBDA} PD={10*LAMBDA+width_N}

* M8 n2 A0 n5 n5 CMOSP W={width_P} L={2*LAMBDA}
* +AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
* +AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

* M9 n2 B0 n5 n5 CMOSP W={width_P} L={2*LAMBDA}
* +AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
* +AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

* M10 n5 Cin vdd vdd CMOSP W={width_P} L={2*LAMBDA}
* +AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
* +AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

* M11 c1 n2 vdd vdd CMOSP W={width_P} L={2*LAMBDA}
* +AS={5*width_P*LAMBDA} PS={10*LAMBDA+width_P}
* +AD={5*width_P*LAMBDA} PD={10*LAMBDA+width_P}

* M12 c1 n2 gnd gnd CMOSN W={width_N} L={2*LAMBDA}
* +AS={5*width_N*LAMBDA} PS={10*LAMBDA+width_N}
* +AD={5*width_N*LAMBDA} PD={10*LAMBDA+width_N}

*CMOSN -> d g s b
*CMOSP -> s g d b

M1 N015 A0 0 N016 CMOSN W={2*width_N} L={2*LAMBDA}
+AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M2 N009 B0 N015 N010 CMOSN W={2*width_N} L={2*LAMBDA}
+AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M3 N004 B0 N009 N005 CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

M4 VDD A0 N004 N001 CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

M5 N009 A0 N014 N011 CMOSN W={2*width_N} L={2*LAMBDA}
+AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M6 N009 B0 N014 N012 CMOSN W={2*width_N} L={2*LAMBDA}
+AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M7 N014 Cin 0 N017 CMOSN W={2*width_N} L={2*LAMBDA}
+AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M8 N003 A0 N009 N006 CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

M9 N003 B0 N009 N007 CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

M10 VDD Cin N003 N002 CMOSP W={2*width_P} L={2*LAMBDA}
+AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P}
+AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}

* .ic v(N009) = 1.8

*Inverter
M11 VDD N009 C1 N008 CMOSP W={width_P} L={2*LAMBDA}
+AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M12 C1 N009 0 N013 CMOSN W={width_N} L={2*LAMBDA}
+AS={5*width_N*LAMBDA} PS={10*LAMBDA+width_N}
+AD={5*width_N*LAMBDA} PD={10*LAMBDA+width_N}


.ends