magic
tech scmos
timestamp 1733209804
<< nwell >>
rect -386 125 -189 178
rect -176 125 -151 178
rect -137 125 -112 178
rect -93 66 -69 118
<< ntransistor >>
rect -82 35 -80 55
rect -371 -207 -369 -187
rect -359 -207 -357 -187
rect -347 -207 -345 -187
rect -335 -207 -333 -187
rect -323 -207 -321 -187
rect -311 -207 -309 -187
rect -299 -207 -297 -187
rect -287 -207 -285 -187
rect -275 -207 -273 -187
rect -263 -207 -261 -187
rect -251 -207 -249 -187
rect -239 -207 -237 -187
rect -227 -207 -225 -187
rect -215 -207 -213 -187
rect -203 -207 -201 -187
rect -165 -207 -163 -187
rect -126 -207 -124 -187
<< ptransistor >>
rect -371 131 -369 171
rect -359 131 -357 171
rect -347 131 -345 171
rect -335 131 -333 171
rect -323 131 -321 171
rect -311 131 -309 171
rect -299 131 -297 171
rect -287 131 -285 171
rect -275 131 -273 171
rect -263 131 -261 171
rect -251 131 -249 171
rect -239 131 -237 171
rect -227 131 -225 171
rect -215 131 -213 171
rect -203 131 -201 171
rect -165 131 -163 171
rect -126 131 -124 171
rect -82 72 -80 112
<< ndiffusion >>
rect -83 35 -82 55
rect -80 35 -79 55
rect -372 -207 -371 -187
rect -369 -207 -368 -187
rect -360 -207 -359 -187
rect -357 -207 -356 -187
rect -348 -207 -347 -187
rect -345 -207 -344 -187
rect -336 -207 -335 -187
rect -333 -207 -332 -187
rect -324 -207 -323 -187
rect -321 -207 -320 -187
rect -312 -207 -311 -187
rect -309 -207 -308 -187
rect -300 -207 -299 -187
rect -297 -207 -296 -187
rect -288 -207 -287 -187
rect -285 -207 -284 -187
rect -276 -207 -275 -187
rect -273 -207 -272 -187
rect -264 -207 -263 -187
rect -261 -207 -260 -187
rect -252 -207 -251 -187
rect -249 -207 -248 -187
rect -240 -207 -239 -187
rect -237 -207 -236 -187
rect -228 -207 -227 -187
rect -225 -207 -224 -187
rect -216 -207 -215 -187
rect -213 -207 -212 -187
rect -204 -207 -203 -187
rect -201 -207 -200 -187
rect -166 -207 -165 -187
rect -163 -207 -162 -187
rect -127 -207 -126 -187
rect -124 -207 -123 -187
<< pdiffusion >>
rect -372 131 -371 171
rect -369 131 -368 171
rect -360 131 -359 171
rect -357 131 -356 171
rect -348 131 -347 171
rect -345 131 -344 171
rect -336 131 -335 171
rect -333 131 -332 171
rect -324 131 -323 171
rect -321 131 -320 171
rect -312 131 -311 171
rect -309 131 -308 171
rect -300 131 -299 171
rect -297 131 -296 171
rect -288 131 -287 171
rect -285 131 -284 171
rect -276 131 -275 171
rect -273 131 -272 171
rect -264 131 -263 171
rect -261 131 -260 171
rect -252 131 -251 171
rect -249 131 -248 171
rect -240 131 -239 171
rect -237 131 -236 171
rect -228 131 -227 171
rect -225 131 -224 171
rect -216 131 -215 171
rect -213 131 -212 171
rect -204 131 -203 171
rect -201 131 -200 171
rect -166 131 -165 171
rect -163 131 -162 171
rect -127 131 -126 171
rect -124 131 -123 171
rect -83 72 -82 112
rect -80 72 -79 112
<< ndcontact >>
rect -87 35 -83 55
rect -79 35 -75 55
rect -376 -207 -372 -187
rect -368 -207 -360 -187
rect -356 -207 -348 -187
rect -344 -207 -336 -187
rect -332 -207 -324 -187
rect -320 -207 -312 -187
rect -308 -207 -300 -187
rect -296 -207 -288 -187
rect -284 -207 -276 -187
rect -272 -207 -264 -187
rect -260 -207 -252 -187
rect -248 -207 -240 -187
rect -236 -207 -228 -187
rect -224 -207 -216 -187
rect -212 -207 -204 -187
rect -200 -207 -196 -187
rect -170 -207 -166 -187
rect -162 -207 -158 -187
rect -131 -207 -127 -187
rect -123 -207 -119 -187
<< pdcontact >>
rect -376 131 -372 171
rect -368 131 -360 171
rect -356 131 -348 171
rect -344 131 -336 171
rect -332 131 -324 171
rect -320 131 -312 171
rect -308 131 -300 171
rect -296 131 -288 171
rect -284 131 -276 171
rect -272 131 -264 171
rect -260 131 -252 171
rect -248 131 -240 171
rect -236 131 -228 171
rect -224 131 -216 171
rect -212 131 -204 171
rect -200 131 -196 171
rect -170 131 -166 171
rect -162 131 -158 171
rect -131 131 -127 171
rect -123 131 -119 171
rect -87 72 -83 112
rect -79 72 -75 112
<< polysilicon >>
rect -371 171 -369 174
rect -359 171 -357 175
rect -347 171 -345 174
rect -335 171 -333 174
rect -323 171 -321 174
rect -311 171 -309 174
rect -299 171 -297 174
rect -287 171 -285 174
rect -275 171 -273 174
rect -263 171 -261 174
rect -251 171 -249 174
rect -239 171 -237 174
rect -227 171 -225 174
rect -215 171 -213 174
rect -203 171 -201 174
rect -165 171 -163 174
rect -126 171 -124 174
rect -371 -187 -369 131
rect -359 -187 -357 131
rect -347 -187 -345 131
rect -335 -187 -333 131
rect -323 -187 -321 131
rect -311 -187 -309 131
rect -299 -187 -297 131
rect -287 -187 -285 131
rect -275 -187 -273 131
rect -263 -187 -261 131
rect -251 -187 -249 131
rect -239 -187 -237 131
rect -227 -187 -225 131
rect -215 -187 -213 131
rect -203 -187 -201 131
rect -165 -187 -163 131
rect -126 -187 -124 131
rect -82 112 -80 118
rect -82 55 -80 72
rect -82 31 -80 35
rect -371 -211 -369 -207
rect -359 -210 -357 -207
rect -347 -210 -345 -207
rect -335 -211 -333 -207
rect -323 -212 -321 -207
rect -311 -212 -309 -207
rect -299 -212 -297 -207
rect -287 -211 -285 -207
rect -275 -211 -273 -207
rect -263 -212 -261 -207
rect -251 -212 -249 -207
rect -239 -212 -237 -207
rect -227 -211 -225 -207
rect -215 -211 -213 -207
rect -203 -211 -201 -207
rect -165 -211 -163 -207
rect -126 -211 -124 -207
<< polycontact >>
rect -376 38 -371 44
rect -364 27 -359 32
rect -345 19 -340 24
rect -340 10 -335 15
rect -328 0 -323 6
rect -316 -9 -311 -4
rect -304 -17 -299 -12
rect -292 -26 -287 -21
rect -280 -35 -275 -30
rect -268 -44 -263 -39
rect -256 -53 -251 -48
rect -244 -62 -239 -57
rect -232 -71 -227 -66
rect -220 -80 -215 -75
rect -208 -89 -203 -84
rect -170 -98 -165 -93
rect -131 -107 -126 -102
rect -87 59 -82 63
<< metal1 >>
rect -386 184 -69 188
rect -376 171 -372 184
rect -318 171 -313 184
rect -234 171 -229 184
rect -354 64 -350 131
rect -342 75 -337 131
rect -294 90 -289 131
rect -282 113 -277 131
rect -270 90 -265 131
rect -259 110 -254 131
rect -222 119 -217 131
rect -211 129 -206 131
rect -200 129 -196 131
rect -169 119 -166 131
rect -222 114 -166 119
rect -162 110 -158 131
rect -259 105 -211 110
rect -206 105 -158 110
rect -294 84 -200 90
rect -342 71 -283 75
rect -130 75 -127 131
rect -276 71 -127 75
rect -123 63 -119 131
rect -87 112 -84 184
rect -79 63 -75 72
rect -349 59 -87 63
rect -79 59 -62 63
rect -354 50 -350 55
rect -415 38 -397 44
rect -387 38 -376 44
rect -415 27 -364 32
rect -376 23 -371 27
rect -376 19 -345 23
rect -340 19 -339 23
rect -376 18 -339 19
rect -414 10 -367 15
rect -361 10 -340 15
rect -416 0 -343 6
rect -337 0 -328 6
rect -413 -9 -380 -4
rect -374 -9 -316 -4
rect -417 -17 -331 -12
rect -326 -17 -304 -12
rect -361 -26 -292 -21
rect -337 -35 -280 -30
rect -326 -44 -268 -39
rect -406 -53 -270 -48
rect -265 -53 -256 -48
rect -410 -62 -258 -57
rect -252 -62 -244 -57
rect -408 -71 -232 -66
rect -252 -80 -220 -75
rect -374 -89 -208 -84
rect -265 -98 -170 -93
rect -398 -107 -397 -102
rect -387 -107 -131 -102
rect -342 -119 -284 -113
rect -354 -187 -350 -182
rect -342 -187 -337 -119
rect -277 -119 -127 -113
rect -294 -132 -200 -127
rect -294 -187 -290 -132
rect -283 -187 -278 -175
rect -270 -187 -266 -132
rect -259 -162 -211 -155
rect -205 -162 -158 -155
rect -259 -187 -255 -162
rect -222 -176 -166 -171
rect -222 -187 -218 -176
rect -200 -187 -196 -186
rect -170 -187 -166 -176
rect -162 -187 -158 -162
rect -131 -187 -127 -119
rect -123 -187 -119 59
rect -79 55 -75 59
rect -376 -217 -372 -207
rect -318 -217 -314 -207
rect -234 -217 -230 -207
rect -87 -217 -83 35
rect -377 -222 -69 -217
<< m2contact >>
rect -283 107 -276 113
rect -211 123 -206 129
rect -200 123 -194 129
rect -211 104 -206 110
rect -200 82 -194 91
rect -283 70 -276 76
rect -355 55 -349 64
rect -397 36 -387 44
rect -367 10 -361 15
rect -343 0 -337 6
rect -380 -9 -374 -4
rect -331 -17 -326 -12
rect -367 -26 -361 -21
rect -343 -35 -337 -29
rect -331 -44 -326 -39
rect -270 -53 -265 -48
rect -258 -62 -252 -57
rect -258 -80 -252 -75
rect -380 -89 -374 -84
rect -270 -98 -265 -93
rect -397 -108 -387 -100
rect -355 -182 -349 -173
rect -284 -120 -277 -112
rect -284 -175 -276 -167
rect -200 -133 -195 -126
rect -211 -162 -205 -155
rect -211 -187 -205 -180
rect -200 -186 -195 -181
<< metal2 >>
rect -211 110 -206 123
rect -282 76 -277 107
rect -200 91 -196 123
rect -396 -100 -388 36
rect -380 -84 -374 -9
rect -367 -21 -361 10
rect -354 -173 -350 55
rect -343 -29 -337 0
rect -331 -39 -326 -17
rect -270 -93 -266 -53
rect -258 -75 -253 -62
rect -283 -167 -278 -120
rect -210 -180 -206 -162
rect -354 -187 -350 -182
rect -200 -181 -196 -133
rect -200 -187 -196 -186
<< labels >>
rlabel metal1 -82 187 -82 187 5 vdd
rlabel metal1 -82 -219 -82 -219 1 gnd
rlabel metal1 -413 39 -408 44 1 a3
rlabel metal1 -412 27 -407 32 1 b3
rlabel metal1 -413 10 -407 15 1 b2
rlabel metal1 -413 1 -407 6 1 a2
rlabel metal1 -412 -9 -407 -4 1 a1
rlabel metal1 -413 -17 -407 -12 1 b1
rlabel metal1 -403 -52 -398 -48 1 b0
rlabel metal1 -402 -62 -397 -58 1 a0
rlabel metal1 -401 -71 -396 -67 1 cin
rlabel metal1 -71 59 -67 63 1 cout_new
<< end >>
