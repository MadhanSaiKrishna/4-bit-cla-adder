magic
tech scmos
timestamp 1733157156
<< nwell >>
rect -420 33 -383 132
rect -370 35 -344 132
rect -324 35 -298 132
rect -292 36 -264 88
<< ntransistor >>
rect -277 5 -275 25
rect -408 -43 -406 -3
rect -357 -40 -355 0
rect -345 -40 -343 0
rect -311 -40 -309 0
rect -299 -40 -297 0
<< ptransistor >>
rect -408 41 -406 121
rect -396 41 -394 121
rect -357 41 -355 121
rect -311 41 -309 121
rect -277 42 -275 82
<< ndiffusion >>
rect -278 5 -277 25
rect -275 5 -274 25
rect -409 -43 -408 -3
rect -406 -43 -405 -3
rect -358 -40 -357 0
rect -355 -40 -354 0
rect -346 -40 -345 0
rect -343 -40 -342 0
rect -312 -40 -311 0
rect -309 -40 -308 0
rect -300 -40 -299 0
rect -297 -40 -296 0
<< pdiffusion >>
rect -409 41 -408 121
rect -406 41 -405 121
rect -397 41 -396 121
rect -394 41 -393 121
rect -358 41 -357 121
rect -355 41 -354 121
rect -312 41 -311 121
rect -309 41 -308 121
rect -278 42 -277 82
rect -275 42 -274 82
<< ndcontact >>
rect -282 5 -278 25
rect -274 5 -270 25
rect -413 -43 -409 -3
rect -405 -43 -401 -3
rect -362 -40 -358 0
rect -354 -40 -346 0
rect -342 -40 -338 0
rect -316 -40 -312 0
rect -308 -40 -300 0
rect -296 -40 -292 0
<< pdcontact >>
rect -413 41 -409 121
rect -405 41 -397 121
rect -393 41 -389 121
rect -362 41 -358 121
rect -354 41 -350 121
rect -316 41 -312 121
rect -308 41 -304 121
rect -282 42 -278 82
rect -274 42 -270 82
<< polysilicon >>
rect -408 121 -406 125
rect -396 121 -394 125
rect -357 121 -355 125
rect -311 121 -309 125
rect -277 82 -275 88
rect -408 -3 -406 41
rect -396 17 -394 41
rect -357 24 -355 41
rect -311 24 -309 41
rect -277 25 -275 42
rect -357 0 -355 11
rect -345 0 -343 12
rect -311 0 -309 11
rect -299 0 -297 12
rect -277 1 -275 5
rect -408 -49 -406 -43
rect -357 -44 -355 -40
rect -345 -43 -343 -40
rect -311 -44 -309 -40
rect -299 -43 -297 -40
<< polycontact >>
rect -414 12 -408 17
rect -282 28 -277 32
rect -394 20 -388 24
rect -359 20 -353 24
rect -313 20 -307 24
rect -358 11 -354 15
rect -346 12 -342 17
rect -312 11 -308 15
rect -300 12 -296 17
<< metal1 >>
rect -420 127 -278 135
rect -413 121 -409 127
rect -362 121 -358 127
rect -316 121 -312 127
rect -282 82 -278 127
rect -393 31 -389 41
rect -405 27 -389 31
rect -354 32 -350 41
rect -367 28 -329 32
rect -308 32 -304 41
rect -274 33 -270 42
rect -321 28 -282 32
rect -274 29 -256 33
rect -419 12 -414 17
rect -405 15 -401 27
rect -388 20 -382 24
rect -332 24 -329 28
rect -274 25 -270 29
rect -377 20 -359 24
rect -353 20 -335 24
rect -332 20 -313 24
rect -307 20 -296 24
rect -346 17 -342 20
rect -405 11 -358 15
rect -339 15 -335 20
rect -300 17 -296 20
rect -339 11 -312 15
rect -405 -3 -401 11
rect -413 -49 -409 -43
rect -342 -49 -338 -40
rect -296 -49 -292 -40
rect -282 -49 -277 5
rect -417 -54 -277 -49
<< m2contact >>
rect -372 28 -367 33
rect -326 28 -321 33
rect -382 20 -377 25
rect -363 0 -358 5
rect -317 0 -312 5
<< metal2 >>
rect -382 6 -377 20
rect -419 2 -377 6
rect -372 5 -367 28
rect -326 5 -321 28
rect -372 0 -363 5
rect -326 0 -317 5
<< labels >>
rlabel metal1 -385 22 -385 22 1 clk
rlabel metal1 -418 15 -418 15 3 a_in
rlabel metal1 -270 30 -268 32 7 a
rlabel metal1 -405 -53 -405 -53 1 gnd
rlabel metal1 -312 132 -312 132 5 vdd
rlabel metal1 -358 132 -358 132 5 vdd
rlabel metal1 -401 133 -401 133 5 vdd
rlabel metal2 -412 4 -412 4 1 clk
<< end >>
