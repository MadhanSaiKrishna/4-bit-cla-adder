magic
tech scmos
timestamp 1733204499
<< nwell >>
rect -193 62 -48 115
rect -35 62 -10 115
rect 4 62 29 115
rect 40 -8 64 44
<< ntransistor >>
rect 51 -39 53 -19
rect -182 -246 -180 -226
rect -170 -246 -168 -226
rect -158 -246 -156 -226
rect -146 -246 -144 -226
rect -134 -246 -132 -226
rect -122 -246 -120 -226
rect -110 -246 -108 -226
rect -98 -246 -96 -226
rect -86 -246 -84 -226
rect -74 -246 -72 -226
rect -62 -246 -60 -226
rect -24 -246 -22 -226
rect 15 -246 17 -226
<< ptransistor >>
rect -182 68 -180 108
rect -170 68 -168 108
rect -158 68 -156 108
rect -146 68 -144 108
rect -134 68 -132 108
rect -122 68 -120 108
rect -110 68 -108 108
rect -98 68 -96 108
rect -86 68 -84 108
rect -74 68 -72 108
rect -62 68 -60 108
rect -24 68 -22 108
rect 15 68 17 108
rect 51 -2 53 38
<< ndiffusion >>
rect 50 -39 51 -19
rect 53 -39 54 -19
rect -183 -246 -182 -226
rect -180 -246 -179 -226
rect -171 -246 -170 -226
rect -168 -246 -167 -226
rect -159 -246 -158 -226
rect -156 -246 -155 -226
rect -147 -246 -146 -226
rect -144 -246 -143 -226
rect -135 -246 -134 -226
rect -132 -246 -131 -226
rect -123 -246 -122 -226
rect -120 -246 -119 -226
rect -111 -246 -110 -226
rect -108 -246 -107 -226
rect -99 -246 -98 -226
rect -96 -246 -95 -226
rect -87 -246 -86 -226
rect -84 -246 -83 -226
rect -75 -246 -74 -226
rect -72 -246 -71 -226
rect -63 -246 -62 -226
rect -60 -246 -59 -226
rect -25 -246 -24 -226
rect -22 -246 -21 -226
rect 14 -246 15 -226
rect 17 -246 18 -226
<< pdiffusion >>
rect -183 68 -182 108
rect -180 68 -179 108
rect -171 68 -170 108
rect -168 68 -167 108
rect -159 68 -158 108
rect -156 68 -155 108
rect -147 68 -146 108
rect -144 68 -143 108
rect -135 68 -134 108
rect -132 68 -131 108
rect -123 68 -122 108
rect -120 68 -119 108
rect -111 68 -110 108
rect -108 68 -107 108
rect -99 68 -98 108
rect -96 68 -95 108
rect -87 68 -86 108
rect -84 68 -83 108
rect -75 68 -74 108
rect -72 68 -71 108
rect -63 68 -62 108
rect -60 68 -59 108
rect -25 68 -24 108
rect -22 68 -21 108
rect 14 68 15 108
rect 17 68 18 108
rect 50 -2 51 38
rect 53 -2 54 38
<< ndcontact >>
rect 46 -39 50 -19
rect 54 -39 58 -19
rect -187 -246 -183 -226
rect -179 -246 -171 -226
rect -167 -246 -159 -226
rect -155 -246 -147 -226
rect -143 -246 -135 -226
rect -131 -246 -123 -226
rect -119 -246 -111 -226
rect -107 -246 -99 -226
rect -95 -246 -87 -226
rect -83 -246 -75 -226
rect -71 -246 -63 -226
rect -59 -246 -55 -226
rect -29 -246 -25 -226
rect -21 -246 -17 -226
rect 10 -246 14 -226
rect 18 -246 22 -226
<< pdcontact >>
rect -187 68 -183 108
rect -179 68 -171 108
rect -167 68 -159 108
rect -155 68 -147 108
rect -143 68 -135 108
rect -131 68 -123 108
rect -119 68 -111 108
rect -107 68 -99 108
rect -95 68 -87 108
rect -83 68 -75 108
rect -71 68 -63 108
rect -59 68 -55 108
rect -29 68 -25 108
rect -21 68 -17 108
rect 10 68 14 108
rect 18 68 22 108
rect 46 -2 50 38
rect 54 -2 58 38
<< polysilicon >>
rect -182 108 -180 111
rect -170 108 -168 111
rect -158 108 -156 111
rect -146 108 -144 111
rect -134 108 -132 111
rect -122 108 -120 111
rect -110 108 -108 111
rect -98 108 -96 111
rect -86 108 -84 111
rect -74 108 -72 111
rect -62 108 -60 111
rect -24 108 -22 111
rect 15 108 17 111
rect -182 -226 -180 68
rect -170 -226 -168 68
rect -158 -226 -156 68
rect -146 -226 -144 68
rect -134 -226 -132 68
rect -122 -226 -120 68
rect -110 -226 -108 68
rect -98 -226 -96 68
rect -86 -226 -84 68
rect -74 -226 -72 68
rect -62 -226 -60 68
rect -24 -226 -22 68
rect 15 -226 17 68
rect 51 38 53 44
rect 51 -19 53 -2
rect 51 -43 53 -39
rect -182 -251 -180 -246
rect -170 -251 -168 -246
rect -158 -251 -156 -246
rect -146 -250 -144 -246
rect -134 -250 -132 -246
rect -122 -251 -120 -246
rect -110 -251 -108 -246
rect -98 -251 -96 -246
rect -86 -250 -84 -246
rect -74 -250 -72 -246
rect -62 -250 -60 -246
rect -24 -250 -22 -246
rect 15 -250 17 -246
<< polycontact >>
rect -186 -27 -182 -23
rect -174 -36 -170 -32
rect -156 -44 -152 -40
rect -150 -52 -146 -48
rect -138 -62 -134 -58
rect -126 -70 -122 -66
rect -114 -78 -110 -74
rect -102 -87 -98 -82
rect -90 -97 -86 -92
rect -78 -109 -74 -104
rect -66 -119 -62 -114
rect -28 -129 -24 -124
rect 11 -138 15 -133
rect 46 -15 51 -11
<< metal1 >>
rect -193 126 64 130
rect -187 108 -183 126
rect -129 108 -125 126
rect -59 108 -55 126
rect -165 -11 -161 68
rect -153 16 -149 68
rect -105 39 -101 68
rect -93 16 -89 68
rect -81 39 -77 68
rect -69 50 -65 68
rect -28 50 -25 68
rect -69 47 -25 50
rect -21 40 -17 68
rect 11 16 14 68
rect -153 12 14 16
rect 18 -11 22 68
rect 46 38 49 126
rect 54 -11 58 -2
rect -160 -15 46 -11
rect 54 -15 71 -11
rect -160 -16 22 -15
rect -204 -27 -193 -23
rect -187 -27 -186 -23
rect -204 -36 -174 -32
rect -187 -40 -183 -36
rect -187 -44 -156 -40
rect -152 -44 -150 -40
rect -203 -52 -178 -48
rect -173 -52 -150 -48
rect -202 -62 -154 -58
rect -148 -62 -138 -58
rect -201 -70 -142 -66
rect -137 -70 -126 -66
rect -203 -78 -130 -74
rect -124 -78 -114 -74
rect -173 -87 -102 -82
rect -148 -97 -90 -92
rect -142 -109 -141 -104
rect -136 -109 -78 -104
rect -205 -119 -66 -114
rect -124 -129 -28 -124
rect -187 -138 11 -133
rect -153 -177 14 -173
rect -165 -226 -161 -183
rect -153 -226 -149 -177
rect -105 -226 -102 -206
rect -92 -226 -88 -177
rect -80 -226 -77 -205
rect -69 -220 -26 -215
rect -69 -226 -66 -220
rect -29 -226 -26 -220
rect -21 -226 -18 -205
rect 10 -226 14 -177
rect 18 -226 22 -16
rect 54 -19 58 -15
rect -187 -267 -183 -246
rect -129 -267 -125 -246
rect -59 -267 -55 -246
rect 46 -267 50 -39
rect -187 -272 64 -267
<< m2contact >>
rect -106 34 -100 39
rect -82 34 -76 39
rect -21 35 -15 40
rect -166 -17 -160 -11
rect -193 -28 -187 -22
rect -178 -53 -173 -47
rect -154 -63 -148 -57
rect -142 -70 -137 -65
rect -130 -79 -124 -73
rect -178 -88 -173 -81
rect -154 -98 -148 -91
rect -141 -109 -136 -104
rect -130 -130 -124 -124
rect -193 -139 -187 -133
rect -166 -183 -161 -178
rect -106 -206 -101 -201
rect -80 -205 -75 -200
rect -21 -205 -16 -200
<< metal2 >>
rect -100 35 -82 39
rect -76 35 -21 39
rect -165 -11 -161 -10
rect -193 -133 -187 -28
rect -178 -81 -174 -53
rect -165 -178 -161 -17
rect -153 -91 -149 -63
rect -137 -70 -136 -66
rect -142 -104 -136 -70
rect -142 -109 -141 -104
rect -129 -124 -125 -79
rect -101 -205 -80 -201
rect -75 -205 -21 -201
<< labels >>
rlabel metal1 51 129 51 129 5 vdd
rlabel metal1 51 -269 51 -269 1 gnd
rlabel metal1 -198 -27 -193 -23 1 a2
rlabel metal1 -197 -36 -192 -32 1 b2
rlabel metal1 -196 -52 -192 -48 1 b1
rlabel metal1 -196 -62 -192 -58 1 a1
rlabel metal1 -195 -70 -191 -66 1 a0
rlabel metal1 -194 -78 -190 -74 1 b0
rlabel metal1 -194 -119 -189 -114 1 cin
rlabel metal1 63 -15 70 -11 7 c3
<< end >>
