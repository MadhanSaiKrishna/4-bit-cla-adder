magic
tech scmos
timestamp 1733170715
<< nwell >>
rect -386 87 -189 140
rect -176 87 -151 140
rect -137 87 -112 140
rect -93 66 -69 118
<< ntransistor >>
rect -82 35 -80 55
rect -371 14 -369 34
rect -359 14 -357 34
rect -347 14 -345 34
rect -335 14 -333 34
rect -323 14 -321 34
rect -311 14 -309 34
rect -299 14 -297 34
rect -287 14 -285 34
rect -275 14 -273 34
rect -263 14 -261 34
rect -251 14 -249 34
rect -239 14 -237 34
rect -227 14 -225 34
rect -215 14 -213 34
rect -203 14 -201 34
rect -165 14 -163 34
rect -126 14 -124 34
<< ptransistor >>
rect -371 93 -369 133
rect -359 93 -357 133
rect -347 93 -345 133
rect -335 93 -333 133
rect -323 93 -321 133
rect -311 93 -309 133
rect -299 93 -297 133
rect -287 93 -285 133
rect -275 93 -273 133
rect -263 93 -261 133
rect -251 93 -249 133
rect -239 93 -237 133
rect -227 93 -225 133
rect -215 93 -213 133
rect -203 93 -201 133
rect -165 93 -163 133
rect -126 93 -124 133
rect -82 72 -80 112
<< ndiffusion >>
rect -83 35 -82 55
rect -80 35 -79 55
rect -372 14 -371 34
rect -369 14 -368 34
rect -360 14 -359 34
rect -357 14 -356 34
rect -348 14 -347 34
rect -345 14 -344 34
rect -336 14 -335 34
rect -333 14 -332 34
rect -324 14 -323 34
rect -321 14 -320 34
rect -312 14 -311 34
rect -309 14 -308 34
rect -300 14 -299 34
rect -297 14 -296 34
rect -288 14 -287 34
rect -285 14 -284 34
rect -276 14 -275 34
rect -273 14 -272 34
rect -264 14 -263 34
rect -261 14 -260 34
rect -252 14 -251 34
rect -249 14 -248 34
rect -240 14 -239 34
rect -237 14 -236 34
rect -228 14 -227 34
rect -225 14 -224 34
rect -216 14 -215 34
rect -213 14 -212 34
rect -204 14 -203 34
rect -201 14 -200 34
rect -166 14 -165 34
rect -163 14 -162 34
rect -127 14 -126 34
rect -124 14 -123 34
<< pdiffusion >>
rect -372 93 -371 133
rect -369 93 -368 133
rect -360 93 -359 133
rect -357 93 -356 133
rect -348 93 -347 133
rect -345 93 -344 133
rect -336 93 -335 133
rect -333 93 -332 133
rect -324 93 -323 133
rect -321 93 -320 133
rect -312 93 -311 133
rect -309 93 -308 133
rect -300 93 -299 133
rect -297 93 -296 133
rect -288 93 -287 133
rect -285 93 -284 133
rect -276 93 -275 133
rect -273 93 -272 133
rect -264 93 -263 133
rect -261 93 -260 133
rect -252 93 -251 133
rect -249 93 -248 133
rect -240 93 -239 133
rect -237 93 -236 133
rect -228 93 -227 133
rect -225 93 -224 133
rect -216 93 -215 133
rect -213 93 -212 133
rect -204 93 -203 133
rect -201 93 -200 133
rect -166 93 -165 133
rect -163 93 -162 133
rect -127 93 -126 133
rect -124 93 -123 133
rect -83 72 -82 112
rect -80 72 -79 112
<< ndcontact >>
rect -87 35 -83 55
rect -79 35 -75 55
rect -376 14 -372 34
rect -368 14 -360 34
rect -356 14 -348 34
rect -344 14 -336 34
rect -332 14 -324 34
rect -320 14 -312 34
rect -308 14 -300 34
rect -296 14 -288 34
rect -284 14 -276 34
rect -272 14 -264 34
rect -260 14 -252 34
rect -248 14 -240 34
rect -236 14 -228 34
rect -224 14 -216 34
rect -212 14 -204 34
rect -200 14 -196 34
rect -170 14 -166 34
rect -162 14 -158 34
rect -131 14 -127 34
rect -123 14 -119 34
<< pdcontact >>
rect -376 93 -372 133
rect -368 93 -360 133
rect -356 93 -348 133
rect -344 93 -336 133
rect -332 93 -324 133
rect -320 93 -312 133
rect -308 93 -300 133
rect -296 93 -288 133
rect -284 93 -276 133
rect -272 93 -264 133
rect -260 93 -252 133
rect -248 93 -240 133
rect -236 93 -228 133
rect -224 93 -216 133
rect -212 93 -204 133
rect -200 93 -196 133
rect -170 93 -166 133
rect -162 93 -158 133
rect -131 93 -127 133
rect -123 93 -119 133
rect -87 72 -83 112
rect -79 72 -75 112
<< polysilicon >>
rect -371 133 -369 136
rect -359 133 -357 137
rect -347 133 -345 136
rect -335 133 -333 136
rect -323 133 -321 136
rect -311 133 -309 136
rect -299 133 -297 136
rect -287 133 -285 136
rect -275 133 -273 136
rect -263 133 -261 136
rect -251 133 -249 136
rect -239 133 -237 136
rect -227 133 -225 136
rect -215 133 -213 136
rect -203 133 -201 136
rect -165 133 -163 136
rect -126 133 -124 136
rect -82 112 -80 118
rect -371 34 -369 93
rect -359 34 -357 93
rect -347 34 -345 93
rect -335 34 -333 93
rect -323 34 -321 93
rect -311 34 -309 93
rect -299 34 -297 93
rect -287 34 -285 93
rect -275 34 -273 93
rect -263 34 -261 93
rect -251 34 -249 93
rect -239 34 -237 93
rect -227 34 -225 93
rect -215 34 -213 93
rect -203 34 -201 93
rect -165 34 -163 93
rect -126 34 -124 93
rect -82 55 -80 72
rect -82 31 -80 35
rect -371 10 -369 14
rect -359 11 -357 14
rect -347 11 -345 14
rect -335 10 -333 14
rect -323 9 -321 14
rect -311 9 -309 14
rect -299 9 -297 14
rect -287 10 -285 14
rect -275 10 -273 14
rect -263 9 -261 14
rect -251 9 -249 14
rect -239 9 -237 14
rect -227 10 -225 14
rect -215 10 -213 14
rect -203 10 -201 14
rect -165 10 -163 14
rect -126 10 -124 14
<< polycontact >>
rect -87 59 -82 63
<< metal1 >>
rect -386 140 -69 144
rect -169 85 -166 93
rect -162 85 -158 93
rect -130 85 -127 93
rect -123 85 -119 93
rect -87 112 -84 140
rect -79 63 -75 72
rect -101 59 -87 63
rect -79 59 -62 63
rect -79 55 -75 59
rect -87 -3 -83 35
rect -377 -8 -69 -3
<< labels >>
rlabel metal1 -82 143 -82 143 5 vdd
rlabel metal1 -82 -5 -82 -5 1 gnd
<< end >>
