magic
tech scmos
timestamp 1733204889
<< nwell >>
rect -193 62 -48 115
rect -35 62 -10 115
rect 4 62 29 115
rect 40 -8 64 44
<< ntransistor >>
rect 51 -39 53 -19
rect -182 -223 -180 -203
rect -170 -223 -168 -203
rect -158 -223 -156 -203
rect -146 -223 -144 -203
rect -134 -223 -132 -203
rect -122 -223 -120 -203
rect -110 -223 -108 -203
rect -98 -223 -96 -203
rect -86 -223 -84 -203
rect -74 -223 -72 -203
rect -62 -223 -60 -203
rect -24 -223 -22 -203
rect 15 -223 17 -203
<< ptransistor >>
rect -182 68 -180 108
rect -170 68 -168 108
rect -158 68 -156 108
rect -146 68 -144 108
rect -134 68 -132 108
rect -122 68 -120 108
rect -110 68 -108 108
rect -98 68 -96 108
rect -86 68 -84 108
rect -74 68 -72 108
rect -62 68 -60 108
rect -24 68 -22 108
rect 15 68 17 108
rect 51 -2 53 38
<< ndiffusion >>
rect 50 -39 51 -19
rect 53 -39 54 -19
rect -183 -223 -182 -203
rect -180 -223 -179 -203
rect -171 -223 -170 -203
rect -168 -223 -167 -203
rect -159 -223 -158 -203
rect -156 -223 -155 -203
rect -147 -223 -146 -203
rect -144 -223 -143 -203
rect -135 -223 -134 -203
rect -132 -223 -131 -203
rect -123 -223 -122 -203
rect -120 -223 -119 -203
rect -111 -223 -110 -203
rect -108 -223 -107 -203
rect -99 -223 -98 -203
rect -96 -223 -95 -203
rect -87 -223 -86 -203
rect -84 -223 -83 -203
rect -75 -223 -74 -203
rect -72 -223 -71 -203
rect -63 -223 -62 -203
rect -60 -223 -59 -203
rect -25 -223 -24 -203
rect -22 -223 -21 -203
rect 14 -223 15 -203
rect 17 -223 18 -203
<< pdiffusion >>
rect -183 68 -182 108
rect -180 68 -179 108
rect -171 68 -170 108
rect -168 68 -167 108
rect -159 68 -158 108
rect -156 68 -155 108
rect -147 68 -146 108
rect -144 68 -143 108
rect -135 68 -134 108
rect -132 68 -131 108
rect -123 68 -122 108
rect -120 68 -119 108
rect -111 68 -110 108
rect -108 68 -107 108
rect -99 68 -98 108
rect -96 68 -95 108
rect -87 68 -86 108
rect -84 68 -83 108
rect -75 68 -74 108
rect -72 68 -71 108
rect -63 68 -62 108
rect -60 68 -59 108
rect -25 68 -24 108
rect -22 68 -21 108
rect 14 68 15 108
rect 17 68 18 108
rect 50 -2 51 38
rect 53 -2 54 38
<< ndcontact >>
rect 46 -39 50 -19
rect 54 -39 58 -19
rect -187 -223 -183 -203
rect -179 -223 -171 -203
rect -167 -223 -159 -203
rect -155 -223 -147 -203
rect -143 -223 -135 -203
rect -131 -223 -123 -203
rect -119 -223 -111 -203
rect -107 -223 -99 -203
rect -95 -223 -87 -203
rect -83 -223 -75 -203
rect -71 -223 -63 -203
rect -59 -223 -55 -203
rect -29 -223 -25 -203
rect -21 -223 -17 -203
rect 10 -223 14 -203
rect 18 -223 22 -203
<< pdcontact >>
rect -187 68 -183 108
rect -179 68 -171 108
rect -167 68 -159 108
rect -155 68 -147 108
rect -143 68 -135 108
rect -131 68 -123 108
rect -119 68 -111 108
rect -107 68 -99 108
rect -95 68 -87 108
rect -83 68 -75 108
rect -71 68 -63 108
rect -59 68 -55 108
rect -29 68 -25 108
rect -21 68 -17 108
rect 10 68 14 108
rect 18 68 22 108
rect 46 -2 50 38
rect 54 -2 58 38
<< polysilicon >>
rect -182 108 -180 111
rect -170 108 -168 111
rect -158 108 -156 111
rect -146 108 -144 111
rect -134 108 -132 111
rect -122 108 -120 111
rect -110 108 -108 111
rect -98 108 -96 111
rect -86 108 -84 111
rect -74 108 -72 111
rect -62 108 -60 111
rect -24 108 -22 111
rect 15 108 17 111
rect -182 -203 -180 68
rect -170 -203 -168 68
rect -158 -203 -156 68
rect -146 -203 -144 68
rect -134 -203 -132 68
rect -122 -203 -120 68
rect -110 -203 -108 68
rect -98 -203 -96 68
rect -86 -203 -84 68
rect -74 -203 -72 68
rect -62 -203 -60 68
rect -24 -203 -22 68
rect 15 -203 17 68
rect 51 38 53 44
rect 51 -19 53 -2
rect 51 -43 53 -39
rect -182 -228 -180 -223
rect -170 -228 -168 -223
rect -158 -228 -156 -223
rect -146 -227 -144 -223
rect -134 -227 -132 -223
rect -122 -228 -120 -223
rect -110 -228 -108 -223
rect -98 -228 -96 -223
rect -86 -227 -84 -223
rect -74 -227 -72 -223
rect -62 -227 -60 -223
rect -24 -227 -22 -223
rect 15 -227 17 -223
<< polycontact >>
rect -186 -27 -182 -23
rect -174 -36 -170 -32
rect -156 -44 -152 -40
rect -150 -52 -146 -48
rect -138 -62 -134 -58
rect -126 -70 -122 -66
rect -114 -78 -110 -74
rect -102 -87 -98 -82
rect -90 -97 -86 -92
rect -78 -109 -74 -104
rect -66 -119 -62 -114
rect -28 -129 -24 -124
rect 11 -138 15 -133
rect 46 -15 51 -11
<< metal1 >>
rect -193 126 64 130
rect -187 108 -183 126
rect -129 108 -125 126
rect -59 108 -55 126
rect -165 -11 -161 68
rect -153 16 -149 68
rect -105 39 -101 68
rect -93 16 -89 68
rect -81 39 -77 68
rect -69 50 -65 68
rect -28 50 -25 68
rect -69 47 -25 50
rect -21 40 -17 68
rect 11 16 14 68
rect -153 12 14 16
rect 18 -11 22 68
rect 46 38 49 126
rect 54 -11 58 -2
rect -160 -15 46 -11
rect 54 -15 71 -11
rect -160 -16 22 -15
rect -204 -27 -193 -23
rect -187 -27 -186 -23
rect -204 -36 -174 -32
rect -187 -40 -183 -36
rect -187 -44 -156 -40
rect -152 -44 -150 -40
rect -203 -52 -178 -48
rect -173 -52 -150 -48
rect -202 -62 -154 -58
rect -148 -62 -138 -58
rect -201 -70 -142 -66
rect -137 -70 -126 -66
rect -203 -78 -130 -74
rect -124 -78 -114 -74
rect -173 -87 -102 -82
rect -148 -97 -90 -92
rect -142 -109 -141 -104
rect -136 -109 -78 -104
rect -205 -119 -66 -114
rect -124 -129 -28 -124
rect -187 -138 11 -133
rect -153 -154 14 -150
rect -165 -203 -161 -160
rect -153 -203 -149 -154
rect -105 -203 -102 -183
rect -92 -203 -88 -154
rect -80 -203 -77 -182
rect -69 -197 -26 -192
rect -69 -203 -66 -197
rect -29 -203 -26 -197
rect -21 -203 -18 -182
rect 10 -203 14 -154
rect 18 -203 22 -16
rect 54 -19 58 -15
rect -187 -244 -183 -223
rect -129 -244 -125 -223
rect -59 -244 -55 -223
rect 46 -244 50 -39
rect -187 -249 64 -244
<< m2contact >>
rect -106 34 -100 39
rect -82 34 -76 39
rect -21 35 -15 40
rect -166 -17 -160 -11
rect -193 -28 -187 -22
rect -178 -53 -173 -47
rect -154 -63 -148 -57
rect -142 -70 -137 -65
rect -130 -79 -124 -73
rect -178 -88 -173 -81
rect -154 -98 -148 -91
rect -141 -109 -136 -104
rect -130 -130 -124 -124
rect -193 -139 -187 -133
rect -166 -160 -161 -155
rect -106 -183 -101 -178
rect -80 -182 -75 -177
rect -21 -182 -16 -177
<< metal2 >>
rect -100 35 -82 39
rect -76 35 -21 39
rect -165 -11 -161 -10
rect -193 -133 -187 -28
rect -178 -81 -174 -53
rect -165 -155 -161 -17
rect -153 -91 -149 -63
rect -137 -70 -136 -66
rect -142 -104 -136 -70
rect -142 -109 -141 -104
rect -129 -124 -125 -79
rect -101 -182 -80 -178
rect -75 -182 -21 -178
<< labels >>
rlabel metal1 51 129 51 129 5 vdd
rlabel metal1 -198 -27 -193 -23 1 a2
rlabel metal1 -197 -36 -192 -32 1 b2
rlabel metal1 -196 -52 -192 -48 1 b1
rlabel metal1 -196 -62 -192 -58 1 a1
rlabel metal1 -195 -70 -191 -66 1 a0
rlabel metal1 -194 -78 -190 -74 1 b0
rlabel metal1 -194 -119 -189 -114 1 cin
rlabel metal1 63 -15 70 -11 7 c3
rlabel metal1 51 -246 51 -246 1 gnd
<< end >>
