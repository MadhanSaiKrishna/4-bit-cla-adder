* SPICE3 file created from two_inp_xor.ext - technology: scmos
.include TSMC_180nm.txt
.option scale=0.09u

.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd
Vdd vdd gnd 'SUPPLY'
V1 a0 gnd pulse 0 1.8 0 10p 10p 200n 400n
V2 b0 gnd pulse 0 1.8 0n 0 0 40n 80n  

M1000 vdd a0 a_78_63# w_65_57# CMOSP w=80 l=2
+  ad=1200 pd=360 as=800 ps=180
M1001 a0_inv a0 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=600 ps=200
M1002 b0_inv b0 vdd w_21_97# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1003 P0 a0_inv a_102_63# w_65_57# CMOSP w=80 l=2
+  ad=800 pd=340 as=800 ps=180
M1004 a0_inv a0 vdd w_n18_n10# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1005 P0 b0 a_90_n42# Gnd CMOSN w=40 l=2
+  ad=400 pd=100 as=400 ps=100
M1006 b0_inv b0 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1007 a_71_n42# a0_inv P0 Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1008 gnd b0_inv a_71_n42# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_90_n42# a0 gnd Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_78_63# b0_inv P0 w_65_57# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_102_63# b0 vdd w_65_57# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0

C0 w_65_57# P0 0.21fF
C1 b0 gnd 0.13fF
C2 b0 a0 0.57fF
C3 a_90_n42# gnd 0.41fF
C4 vdd w_65_57# 0.09fF
C5 a_78_63# P0 0.82fF
C6 a_71_n42# gnd 0.52fF
C7 b0 b0_inv 0.13fF
C8 w_n18_n10# vdd 0.06fF
C9 a0 a_71_n42# 0.09fF
C10 a0_inv b0 0.56fF
C11 a_78_63# vdd 0.88fF
C12 b0_inv w_21_97# 0.06fF
C13 b0_inv a_71_n42# 0.09fF
C14 a_78_63# w_65_57# 0.02fF
C15 a0_inv a_71_n42# 0.43fF
C16 b0 P0 0.09fF
C17 a_90_n42# P0 0.41fF
C18 b0 vdd 0.19fF
C19 a_71_n42# P0 1.02fF
C20 a0 gnd 0.13fF
C21 b0 w_65_57# 0.07fF
C22 w_21_97# vdd 0.08fF
C23 b0_inv gnd 0.21fF
C24 b0_inv a0 0.40fF
C25 a0_inv gnd 0.33fF
C26 a0_inv a0 0.20fF
C27 a0_inv b0_inv 0.08fF
C28 a0 P0 0.09fF
C29 a_102_63# P0 0.82fF
C30 a0 vdd 0.09fF
C31 b0_inv P0 0.12fF
C32 a0_inv P0 0.09fF
C33 vdd a_102_63# 0.88fF
C34 b0 w_21_97# 0.08fF
C35 a0 w_65_57# 0.07fF
C36 b0 a_71_n42# 0.09fF
C37 b0_inv vdd 0.44fF
C38 a0_inv vdd 0.41fF
C39 a_90_n42# a_71_n42# 0.08fF
C40 w_n18_n10# a0 0.24fF
C41 w_65_57# a_102_63# 0.02fF
C42 b0_inv w_65_57# 0.07fF
C43 a0_inv w_65_57# 0.07fF
C44 w_n18_n10# a0_inv 0.06fF
C45 vdd P0 0.05fF
C46 a_90_n42# Gnd 0.02fF
C47 a_71_n42# Gnd 0.26fF
C48 a_102_63# Gnd 0.00fF
C49 a_78_63# Gnd 0.00fF
C50 P0 Gnd 0.64fF
C51 gnd Gnd 0.57fF
C52 vdd Gnd 0.01fF
C53 a0_inv Gnd 0.70fF
C54 a0 Gnd 0.17fF
C55 b0_inv Gnd 0.76fF
C56 b0 Gnd 0.51fF
C57 w_n18_n10# Gnd 1.25fF
C58 w_65_57# Gnd 5.54fF
C59 w_21_97# Gnd 1.25fF

.tran 0.1n 1u

.control
set hcopypscolor = 1 
set color0=white
set color1=black
run

plot V(a0) V(b0)+2 V(p0)+4

.endc
.end