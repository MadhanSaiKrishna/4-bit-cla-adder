magic
tech scmos
timestamp 1733225263
<< nwell >>
rect 692 883 889 936
rect 902 883 927 936
rect 941 883 966 936
rect 985 824 1009 876
rect 686 449 831 502
rect 844 449 869 502
rect 883 449 908 502
rect 919 379 943 431
rect -189 88 -152 187
rect -139 90 -113 187
rect -93 90 -67 187
rect -61 91 -33 143
rect -21 88 16 187
rect 29 90 55 187
rect 75 90 101 187
rect 107 91 135 143
rect 145 88 182 187
rect 195 90 221 187
rect 241 90 267 187
rect 273 91 301 143
rect 310 88 347 187
rect 360 90 386 187
rect 406 90 432 187
rect 438 91 466 143
rect 693 44 801 96
rect 815 44 839 96
rect 870 16 894 68
rect -190 -163 -153 -64
rect -140 -161 -114 -64
rect -94 -161 -68 -64
rect -62 -160 -34 -108
rect -22 -163 15 -64
rect 28 -161 54 -64
rect 74 -161 100 -64
rect 106 -160 134 -108
rect 144 -163 181 -64
rect 194 -161 220 -64
rect 240 -161 266 -64
rect 272 -160 300 -108
rect 309 -163 346 -64
rect 359 -161 385 -64
rect 405 -161 431 -64
rect 437 -160 465 -108
rect 677 -314 743 -261
rect 749 -314 775 -261
rect 782 -313 806 -261
<< ntransistor >>
rect 996 793 998 813
rect 707 551 709 571
rect 719 551 721 571
rect 731 551 733 571
rect 743 551 745 571
rect 755 551 757 571
rect 767 551 769 571
rect 779 551 781 571
rect 791 551 793 571
rect 803 551 805 571
rect 815 551 817 571
rect 827 551 829 571
rect 839 551 841 571
rect 851 551 853 571
rect 863 551 865 571
rect 875 551 877 571
rect 913 551 915 571
rect 952 551 954 571
rect 930 348 932 368
rect -46 60 -44 80
rect -177 12 -175 52
rect -126 15 -124 55
rect -114 15 -112 55
rect -80 15 -78 55
rect -68 15 -66 55
rect 122 60 124 80
rect -9 12 -7 52
rect 42 15 44 55
rect 54 15 56 55
rect 88 15 90 55
rect 100 15 102 55
rect 697 164 699 184
rect 709 164 711 184
rect 721 164 723 184
rect 733 164 735 184
rect 745 164 747 184
rect 757 164 759 184
rect 769 164 771 184
rect 781 164 783 184
rect 793 164 795 184
rect 805 164 807 184
rect 817 164 819 184
rect 855 164 857 184
rect 894 164 896 184
rect 288 60 290 80
rect 157 12 159 52
rect 208 15 210 55
rect 220 15 222 55
rect 254 15 256 55
rect 266 15 268 55
rect 453 60 455 80
rect 322 12 324 52
rect 373 15 375 55
rect 385 15 387 55
rect 419 15 421 55
rect 431 15 433 55
rect -47 -191 -45 -171
rect -178 -239 -176 -199
rect -127 -236 -125 -196
rect -115 -236 -113 -196
rect -81 -236 -79 -196
rect -69 -236 -67 -196
rect 121 -191 123 -171
rect -10 -239 -8 -199
rect 41 -236 43 -196
rect 53 -236 55 -196
rect 87 -236 89 -196
rect 99 -236 101 -196
rect 881 -15 883 5
rect 704 -123 706 -103
rect 716 -123 718 -103
rect 728 -123 730 -103
rect 740 -123 742 -103
rect 752 -123 754 -103
rect 764 -123 766 -103
rect 776 -123 778 -103
rect 788 -123 790 -103
rect 826 -111 828 -91
rect 287 -191 289 -171
rect 156 -239 158 -199
rect 207 -236 209 -196
rect 219 -236 221 -196
rect 253 -236 255 -196
rect 265 -236 267 -196
rect 452 -191 454 -171
rect 321 -239 323 -199
rect 372 -236 374 -196
rect 384 -236 386 -196
rect 418 -236 420 -196
rect 430 -236 432 -196
rect 688 -370 690 -350
rect 700 -370 702 -350
rect 712 -370 714 -350
rect 724 -370 726 -350
rect 761 -370 763 -350
rect 793 -393 795 -373
<< ptransistor >>
rect 707 889 709 929
rect 719 889 721 929
rect 731 889 733 929
rect 743 889 745 929
rect 755 889 757 929
rect 767 889 769 929
rect 779 889 781 929
rect 791 889 793 929
rect 803 889 805 929
rect 815 889 817 929
rect 827 889 829 929
rect 839 889 841 929
rect 851 889 853 929
rect 863 889 865 929
rect 875 889 877 929
rect 913 889 915 929
rect 952 889 954 929
rect 996 830 998 870
rect 697 455 699 495
rect 709 455 711 495
rect 721 455 723 495
rect 733 455 735 495
rect 745 455 747 495
rect 757 455 759 495
rect 769 455 771 495
rect 781 455 783 495
rect 793 455 795 495
rect 805 455 807 495
rect 817 455 819 495
rect 855 455 857 495
rect 894 455 896 495
rect 930 385 932 425
rect -177 96 -175 176
rect -165 96 -163 176
rect -126 96 -124 176
rect -80 96 -78 176
rect -46 97 -44 137
rect -9 96 -7 176
rect 3 96 5 176
rect 42 96 44 176
rect 88 96 90 176
rect 122 97 124 137
rect 157 96 159 176
rect 169 96 171 176
rect 208 96 210 176
rect 254 96 256 176
rect 288 97 290 137
rect 322 96 324 176
rect 334 96 336 176
rect 373 96 375 176
rect 419 96 421 176
rect 453 97 455 137
rect 704 50 706 90
rect 716 50 718 90
rect 728 50 730 90
rect 740 50 742 90
rect 752 50 754 90
rect 764 50 766 90
rect 776 50 778 90
rect 788 50 790 90
rect 826 50 828 90
rect -178 -155 -176 -75
rect -166 -155 -164 -75
rect -127 -155 -125 -75
rect -81 -155 -79 -75
rect -47 -154 -45 -114
rect -10 -155 -8 -75
rect 2 -155 4 -75
rect 41 -155 43 -75
rect 87 -155 89 -75
rect 121 -154 123 -114
rect 156 -155 158 -75
rect 168 -155 170 -75
rect 207 -155 209 -75
rect 253 -155 255 -75
rect 287 -154 289 -114
rect 321 -155 323 -75
rect 333 -155 335 -75
rect 372 -155 374 -75
rect 418 -155 420 -75
rect 881 22 883 62
rect 452 -154 454 -114
rect 688 -308 690 -268
rect 700 -308 702 -268
rect 712 -308 714 -268
rect 724 -308 726 -268
rect 761 -308 763 -268
rect 793 -307 795 -267
<< ndiffusion >>
rect 995 793 996 813
rect 998 793 999 813
rect 706 551 707 571
rect 709 551 710 571
rect 718 551 719 571
rect 721 551 722 571
rect 730 551 731 571
rect 733 551 734 571
rect 742 551 743 571
rect 745 551 746 571
rect 754 551 755 571
rect 757 551 758 571
rect 766 551 767 571
rect 769 551 770 571
rect 778 551 779 571
rect 781 551 782 571
rect 790 551 791 571
rect 793 551 794 571
rect 802 551 803 571
rect 805 551 806 571
rect 814 551 815 571
rect 817 551 818 571
rect 826 551 827 571
rect 829 551 830 571
rect 838 551 839 571
rect 841 551 842 571
rect 850 551 851 571
rect 853 551 854 571
rect 862 551 863 571
rect 865 551 866 571
rect 874 551 875 571
rect 877 551 878 571
rect 912 551 913 571
rect 915 551 916 571
rect 951 551 952 571
rect 954 551 955 571
rect 929 348 930 368
rect 932 348 933 368
rect -47 60 -46 80
rect -44 60 -43 80
rect -178 12 -177 52
rect -175 12 -174 52
rect -127 15 -126 55
rect -124 15 -123 55
rect -115 15 -114 55
rect -112 15 -111 55
rect -81 15 -80 55
rect -78 15 -77 55
rect -69 15 -68 55
rect -66 15 -65 55
rect 121 60 122 80
rect 124 60 125 80
rect -10 12 -9 52
rect -7 12 -6 52
rect 41 15 42 55
rect 44 15 45 55
rect 53 15 54 55
rect 56 15 57 55
rect 87 15 88 55
rect 90 15 91 55
rect 99 15 100 55
rect 102 15 103 55
rect 696 164 697 184
rect 699 164 700 184
rect 708 164 709 184
rect 711 164 712 184
rect 720 164 721 184
rect 723 164 724 184
rect 732 164 733 184
rect 735 164 736 184
rect 744 164 745 184
rect 747 164 748 184
rect 756 164 757 184
rect 759 164 760 184
rect 768 164 769 184
rect 771 164 772 184
rect 780 164 781 184
rect 783 164 784 184
rect 792 164 793 184
rect 795 164 796 184
rect 804 164 805 184
rect 807 164 808 184
rect 816 164 817 184
rect 819 164 820 184
rect 854 164 855 184
rect 857 164 858 184
rect 893 164 894 184
rect 896 164 897 184
rect 287 60 288 80
rect 290 60 291 80
rect 156 12 157 52
rect 159 12 160 52
rect 207 15 208 55
rect 210 15 211 55
rect 219 15 220 55
rect 222 15 223 55
rect 253 15 254 55
rect 256 15 257 55
rect 265 15 266 55
rect 268 15 269 55
rect 452 60 453 80
rect 455 60 456 80
rect 321 12 322 52
rect 324 12 325 52
rect 372 15 373 55
rect 375 15 376 55
rect 384 15 385 55
rect 387 15 388 55
rect 418 15 419 55
rect 421 15 422 55
rect 430 15 431 55
rect 433 15 434 55
rect -48 -191 -47 -171
rect -45 -191 -44 -171
rect -179 -239 -178 -199
rect -176 -239 -175 -199
rect -128 -236 -127 -196
rect -125 -236 -124 -196
rect -116 -236 -115 -196
rect -113 -236 -112 -196
rect -82 -236 -81 -196
rect -79 -236 -78 -196
rect -70 -236 -69 -196
rect -67 -236 -66 -196
rect 120 -191 121 -171
rect 123 -191 124 -171
rect -11 -239 -10 -199
rect -8 -239 -7 -199
rect 40 -236 41 -196
rect 43 -236 44 -196
rect 52 -236 53 -196
rect 55 -236 56 -196
rect 86 -236 87 -196
rect 89 -236 90 -196
rect 98 -236 99 -196
rect 101 -236 102 -196
rect 880 -15 881 5
rect 883 -15 884 5
rect 703 -123 704 -103
rect 706 -123 707 -103
rect 715 -123 716 -103
rect 718 -123 719 -103
rect 727 -123 728 -103
rect 730 -123 731 -103
rect 739 -123 740 -103
rect 742 -123 743 -103
rect 751 -123 752 -103
rect 754 -123 755 -103
rect 763 -123 764 -103
rect 766 -123 767 -103
rect 775 -123 776 -103
rect 778 -123 779 -103
rect 787 -123 788 -103
rect 790 -123 791 -103
rect 825 -111 826 -91
rect 828 -111 829 -91
rect 286 -191 287 -171
rect 289 -191 290 -171
rect 155 -239 156 -199
rect 158 -239 159 -199
rect 206 -236 207 -196
rect 209 -236 210 -196
rect 218 -236 219 -196
rect 221 -236 222 -196
rect 252 -236 253 -196
rect 255 -236 256 -196
rect 264 -236 265 -196
rect 267 -236 268 -196
rect 451 -191 452 -171
rect 454 -191 455 -171
rect 320 -239 321 -199
rect 323 -239 324 -199
rect 371 -236 372 -196
rect 374 -236 375 -196
rect 383 -236 384 -196
rect 386 -236 387 -196
rect 417 -236 418 -196
rect 420 -236 421 -196
rect 429 -236 430 -196
rect 432 -236 433 -196
rect 687 -370 688 -350
rect 690 -370 691 -350
rect 699 -370 700 -350
rect 702 -370 703 -350
rect 711 -370 712 -350
rect 714 -370 715 -350
rect 723 -370 724 -350
rect 726 -370 727 -350
rect 760 -370 761 -350
rect 763 -370 764 -350
rect 792 -393 793 -373
rect 795 -393 796 -373
<< pdiffusion >>
rect 706 889 707 929
rect 709 889 710 929
rect 718 889 719 929
rect 721 889 722 929
rect 730 889 731 929
rect 733 889 734 929
rect 742 889 743 929
rect 745 889 746 929
rect 754 889 755 929
rect 757 889 758 929
rect 766 889 767 929
rect 769 889 770 929
rect 778 889 779 929
rect 781 889 782 929
rect 790 889 791 929
rect 793 889 794 929
rect 802 889 803 929
rect 805 889 806 929
rect 814 889 815 929
rect 817 889 818 929
rect 826 889 827 929
rect 829 889 830 929
rect 838 889 839 929
rect 841 889 842 929
rect 850 889 851 929
rect 853 889 854 929
rect 862 889 863 929
rect 865 889 866 929
rect 874 889 875 929
rect 877 889 878 929
rect 912 889 913 929
rect 915 889 916 929
rect 951 889 952 929
rect 954 889 955 929
rect 995 830 996 870
rect 998 830 999 870
rect 696 455 697 495
rect 699 455 700 495
rect 708 455 709 495
rect 711 455 712 495
rect 720 455 721 495
rect 723 455 724 495
rect 732 455 733 495
rect 735 455 736 495
rect 744 455 745 495
rect 747 455 748 495
rect 756 455 757 495
rect 759 455 760 495
rect 768 455 769 495
rect 771 455 772 495
rect 780 455 781 495
rect 783 455 784 495
rect 792 455 793 495
rect 795 455 796 495
rect 804 455 805 495
rect 807 455 808 495
rect 816 455 817 495
rect 819 455 820 495
rect 854 455 855 495
rect 857 455 858 495
rect 893 455 894 495
rect 896 455 897 495
rect 929 385 930 425
rect 932 385 933 425
rect -178 96 -177 176
rect -175 96 -174 176
rect -166 96 -165 176
rect -163 96 -162 176
rect -127 96 -126 176
rect -124 96 -123 176
rect -81 96 -80 176
rect -78 96 -77 176
rect -47 97 -46 137
rect -44 97 -43 137
rect -10 96 -9 176
rect -7 96 -6 176
rect 2 96 3 176
rect 5 96 6 176
rect 41 96 42 176
rect 44 96 45 176
rect 87 96 88 176
rect 90 96 91 176
rect 121 97 122 137
rect 124 97 125 137
rect 156 96 157 176
rect 159 96 160 176
rect 168 96 169 176
rect 171 96 172 176
rect 207 96 208 176
rect 210 96 211 176
rect 253 96 254 176
rect 256 96 257 176
rect 287 97 288 137
rect 290 97 291 137
rect 321 96 322 176
rect 324 96 325 176
rect 333 96 334 176
rect 336 96 337 176
rect 372 96 373 176
rect 375 96 376 176
rect 418 96 419 176
rect 421 96 422 176
rect 452 97 453 137
rect 455 97 456 137
rect 703 50 704 90
rect 706 50 707 90
rect 715 50 716 90
rect 718 50 719 90
rect 727 50 728 90
rect 730 50 731 90
rect 739 50 740 90
rect 742 50 743 90
rect 751 50 752 90
rect 754 50 755 90
rect 763 50 764 90
rect 766 50 767 90
rect 775 50 776 90
rect 778 50 779 90
rect 787 50 788 90
rect 790 50 791 90
rect 825 50 826 90
rect 828 50 829 90
rect -179 -155 -178 -75
rect -176 -155 -175 -75
rect -167 -155 -166 -75
rect -164 -155 -163 -75
rect -128 -155 -127 -75
rect -125 -155 -124 -75
rect -82 -155 -81 -75
rect -79 -155 -78 -75
rect -48 -154 -47 -114
rect -45 -154 -44 -114
rect -11 -155 -10 -75
rect -8 -155 -7 -75
rect 1 -155 2 -75
rect 4 -155 5 -75
rect 40 -155 41 -75
rect 43 -155 44 -75
rect 86 -155 87 -75
rect 89 -155 90 -75
rect 120 -154 121 -114
rect 123 -154 124 -114
rect 155 -155 156 -75
rect 158 -155 159 -75
rect 167 -155 168 -75
rect 170 -155 171 -75
rect 206 -155 207 -75
rect 209 -155 210 -75
rect 252 -155 253 -75
rect 255 -155 256 -75
rect 286 -154 287 -114
rect 289 -154 290 -114
rect 320 -155 321 -75
rect 323 -155 324 -75
rect 332 -155 333 -75
rect 335 -155 336 -75
rect 371 -155 372 -75
rect 374 -155 375 -75
rect 417 -155 418 -75
rect 420 -155 421 -75
rect 880 22 881 62
rect 883 22 884 62
rect 451 -154 452 -114
rect 454 -154 455 -114
rect 687 -308 688 -268
rect 690 -308 691 -268
rect 699 -308 700 -268
rect 702 -308 703 -268
rect 711 -308 712 -268
rect 714 -308 715 -268
rect 723 -308 724 -268
rect 726 -308 727 -268
rect 760 -308 761 -268
rect 763 -308 764 -268
rect 792 -307 793 -267
rect 795 -307 796 -267
<< ndcontact >>
rect 991 793 995 813
rect 999 793 1003 813
rect 702 551 706 571
rect 710 551 718 571
rect 722 551 730 571
rect 734 551 742 571
rect 746 551 754 571
rect 758 551 766 571
rect 770 551 778 571
rect 782 551 790 571
rect 794 551 802 571
rect 806 551 814 571
rect 818 551 826 571
rect 830 551 838 571
rect 842 551 850 571
rect 854 551 862 571
rect 866 551 874 571
rect 878 551 882 571
rect 908 551 912 571
rect 916 551 920 571
rect 947 551 951 571
rect 955 551 959 571
rect 925 348 929 368
rect 933 348 937 368
rect -51 60 -47 80
rect -43 60 -39 80
rect -182 12 -178 52
rect -174 12 -170 52
rect -131 15 -127 55
rect -123 15 -115 55
rect -111 15 -107 55
rect -85 15 -81 55
rect -77 15 -69 55
rect -65 15 -61 55
rect 117 60 121 80
rect 125 60 129 80
rect -14 12 -10 52
rect -6 12 -2 52
rect 37 15 41 55
rect 45 15 53 55
rect 57 15 61 55
rect 83 15 87 55
rect 91 15 99 55
rect 103 15 107 55
rect 692 164 696 184
rect 700 164 708 184
rect 712 164 720 184
rect 724 164 732 184
rect 736 164 744 184
rect 748 164 756 184
rect 760 164 768 184
rect 772 164 780 184
rect 784 164 792 184
rect 796 164 804 184
rect 808 164 816 184
rect 820 164 824 184
rect 850 164 854 184
rect 858 164 862 184
rect 889 164 893 184
rect 897 164 901 184
rect 283 60 287 80
rect 291 60 295 80
rect 152 12 156 52
rect 160 12 164 52
rect 203 15 207 55
rect 211 15 219 55
rect 223 15 227 55
rect 249 15 253 55
rect 257 15 265 55
rect 269 15 273 55
rect 448 60 452 80
rect 456 60 460 80
rect 317 12 321 52
rect 325 12 329 52
rect 368 15 372 55
rect 376 15 384 55
rect 388 15 392 55
rect 414 15 418 55
rect 422 15 430 55
rect 434 15 438 55
rect -52 -191 -48 -171
rect -44 -191 -40 -171
rect -183 -239 -179 -199
rect -175 -239 -171 -199
rect -132 -236 -128 -196
rect -124 -236 -116 -196
rect -112 -236 -108 -196
rect -86 -236 -82 -196
rect -78 -236 -70 -196
rect -66 -236 -62 -196
rect 116 -191 120 -171
rect 124 -191 128 -171
rect -15 -239 -11 -199
rect -7 -239 -3 -199
rect 36 -236 40 -196
rect 44 -236 52 -196
rect 56 -236 60 -196
rect 82 -236 86 -196
rect 90 -236 98 -196
rect 102 -236 106 -196
rect 876 -15 880 5
rect 884 -15 888 5
rect 699 -123 703 -103
rect 707 -123 715 -103
rect 719 -123 727 -103
rect 731 -123 739 -103
rect 743 -123 751 -103
rect 755 -123 763 -103
rect 767 -123 775 -103
rect 779 -123 787 -103
rect 791 -123 795 -103
rect 821 -111 825 -91
rect 829 -111 833 -91
rect 282 -191 286 -171
rect 290 -191 294 -171
rect 151 -239 155 -199
rect 159 -239 163 -199
rect 202 -236 206 -196
rect 210 -236 218 -196
rect 222 -236 226 -196
rect 248 -236 252 -196
rect 256 -236 264 -196
rect 268 -236 272 -196
rect 447 -191 451 -171
rect 455 -191 459 -171
rect 316 -239 320 -199
rect 324 -239 328 -199
rect 367 -236 371 -196
rect 375 -236 383 -196
rect 387 -236 391 -196
rect 413 -236 417 -196
rect 421 -236 429 -196
rect 433 -236 437 -196
rect 683 -370 687 -350
rect 691 -370 699 -350
rect 703 -370 711 -350
rect 715 -370 723 -350
rect 727 -370 731 -350
rect 756 -370 760 -350
rect 764 -370 768 -350
rect 788 -393 792 -373
rect 796 -393 800 -373
<< pdcontact >>
rect 702 889 706 929
rect 710 889 718 929
rect 722 889 730 929
rect 734 889 742 929
rect 746 889 754 929
rect 758 889 766 929
rect 770 889 778 929
rect 782 889 790 929
rect 794 889 802 929
rect 806 889 814 929
rect 818 889 826 929
rect 830 889 838 929
rect 842 889 850 929
rect 854 889 862 929
rect 866 889 874 929
rect 878 889 882 929
rect 908 889 912 929
rect 916 889 920 929
rect 947 889 951 929
rect 955 889 959 929
rect 991 830 995 870
rect 999 830 1003 870
rect 692 455 696 495
rect 700 455 708 495
rect 712 455 720 495
rect 724 455 732 495
rect 736 455 744 495
rect 748 455 756 495
rect 760 455 768 495
rect 772 455 780 495
rect 784 455 792 495
rect 796 455 804 495
rect 808 455 816 495
rect 820 455 824 495
rect 850 455 854 495
rect 858 455 862 495
rect 889 455 893 495
rect 897 455 901 495
rect 925 385 929 425
rect 933 385 937 425
rect -182 96 -178 176
rect -174 96 -166 176
rect -162 96 -158 176
rect -131 96 -127 176
rect -123 96 -119 176
rect -85 96 -81 176
rect -77 96 -73 176
rect -51 97 -47 137
rect -43 97 -39 137
rect -14 96 -10 176
rect -6 96 2 176
rect 6 96 10 176
rect 37 96 41 176
rect 45 96 49 176
rect 83 96 87 176
rect 91 96 95 176
rect 117 97 121 137
rect 125 97 129 137
rect 152 96 156 176
rect 160 96 168 176
rect 172 96 176 176
rect 203 96 207 176
rect 211 96 215 176
rect 249 96 253 176
rect 257 96 261 176
rect 283 97 287 137
rect 291 97 295 137
rect 317 96 321 176
rect 325 96 333 176
rect 337 96 341 176
rect 368 96 372 176
rect 376 96 380 176
rect 414 96 418 176
rect 422 96 426 176
rect 448 97 452 137
rect 456 97 460 137
rect 699 50 703 90
rect 707 50 715 90
rect 719 50 727 90
rect 731 50 739 90
rect 743 50 751 90
rect 755 50 763 90
rect 767 50 775 90
rect 779 50 787 90
rect 791 50 795 90
rect 821 50 825 90
rect 829 50 833 90
rect -183 -155 -179 -75
rect -175 -155 -167 -75
rect -163 -155 -159 -75
rect -132 -155 -128 -75
rect -124 -155 -120 -75
rect -86 -155 -82 -75
rect -78 -155 -74 -75
rect -52 -154 -48 -114
rect -44 -154 -40 -114
rect -15 -155 -11 -75
rect -7 -155 1 -75
rect 5 -155 9 -75
rect 36 -155 40 -75
rect 44 -155 48 -75
rect 82 -155 86 -75
rect 90 -155 94 -75
rect 116 -154 120 -114
rect 124 -154 128 -114
rect 151 -155 155 -75
rect 159 -155 167 -75
rect 171 -155 175 -75
rect 202 -155 206 -75
rect 210 -155 214 -75
rect 248 -155 252 -75
rect 256 -155 260 -75
rect 282 -154 286 -114
rect 290 -154 294 -114
rect 316 -155 320 -75
rect 324 -155 332 -75
rect 336 -155 340 -75
rect 367 -155 371 -75
rect 375 -155 379 -75
rect 413 -155 417 -75
rect 421 -155 425 -75
rect 876 22 880 62
rect 884 22 888 62
rect 447 -154 451 -114
rect 455 -154 459 -114
rect 683 -308 687 -268
rect 691 -308 699 -268
rect 703 -308 711 -268
rect 715 -308 723 -268
rect 727 -308 731 -268
rect 756 -308 760 -268
rect 764 -308 768 -268
rect 788 -307 792 -267
rect 796 -307 800 -267
<< polysilicon >>
rect 707 929 709 932
rect 719 929 721 933
rect 731 929 733 932
rect 743 929 745 932
rect 755 929 757 932
rect 767 929 769 932
rect 779 929 781 932
rect 791 929 793 932
rect 803 929 805 932
rect 815 929 817 932
rect 827 929 829 932
rect 839 929 841 932
rect 851 929 853 932
rect 863 929 865 932
rect 875 929 877 932
rect 913 929 915 932
rect 952 929 954 932
rect 707 571 709 889
rect 719 571 721 889
rect 731 571 733 889
rect 743 571 745 889
rect 755 571 757 889
rect 767 571 769 889
rect 779 571 781 889
rect 791 571 793 889
rect 803 571 805 889
rect 815 571 817 889
rect 827 571 829 889
rect 839 571 841 889
rect 851 571 853 889
rect 863 571 865 889
rect 875 571 877 889
rect 913 571 915 889
rect 952 571 954 889
rect 996 870 998 876
rect 996 813 998 830
rect 996 789 998 793
rect 707 547 709 551
rect 719 548 721 551
rect 731 548 733 551
rect 743 547 745 551
rect 755 546 757 551
rect 767 546 769 551
rect 779 546 781 551
rect 791 547 793 551
rect 803 547 805 551
rect 815 546 817 551
rect 827 546 829 551
rect 839 546 841 551
rect 851 547 853 551
rect 863 547 865 551
rect 875 547 877 551
rect 913 547 915 551
rect 952 547 954 551
rect 697 495 699 498
rect 709 495 711 498
rect 721 495 723 498
rect 733 495 735 498
rect 745 495 747 498
rect 757 495 759 498
rect 769 495 771 498
rect 781 495 783 498
rect 793 495 795 498
rect 805 495 807 498
rect 817 495 819 498
rect 855 495 857 498
rect 894 495 896 498
rect 697 184 699 455
rect 709 184 711 455
rect 721 184 723 455
rect 733 184 735 455
rect 745 184 747 455
rect 757 184 759 455
rect 769 184 771 455
rect 781 184 783 455
rect 793 184 795 455
rect 805 184 807 455
rect 817 184 819 455
rect 855 184 857 455
rect 894 184 896 455
rect 930 425 932 431
rect 930 368 932 385
rect 930 344 932 348
rect -177 176 -175 180
rect -165 176 -163 180
rect -126 176 -124 180
rect -80 176 -78 180
rect -9 176 -7 180
rect 3 176 5 180
rect 42 176 44 180
rect 88 176 90 180
rect 157 176 159 180
rect 169 176 171 180
rect 208 176 210 180
rect 254 176 256 180
rect 322 176 324 180
rect 334 176 336 180
rect 373 176 375 180
rect 419 176 421 180
rect -46 137 -44 143
rect -177 52 -175 96
rect -165 72 -163 96
rect -126 79 -124 96
rect -80 79 -78 96
rect -46 80 -44 97
rect 122 137 124 143
rect -126 55 -124 66
rect -114 55 -112 67
rect -80 55 -78 66
rect -68 55 -66 67
rect -46 56 -44 60
rect -9 52 -7 96
rect 3 72 5 96
rect 42 79 44 96
rect 88 79 90 96
rect 122 80 124 97
rect 288 137 290 143
rect 42 55 44 66
rect 54 55 56 67
rect 88 55 90 66
rect 100 55 102 67
rect 122 56 124 60
rect -177 6 -175 12
rect -126 11 -124 15
rect -114 12 -112 15
rect -80 11 -78 15
rect -68 12 -66 15
rect 157 52 159 96
rect 169 72 171 96
rect 208 79 210 96
rect 254 79 256 96
rect 288 80 290 97
rect 697 159 699 164
rect 709 159 711 164
rect 721 159 723 164
rect 733 160 735 164
rect 745 160 747 164
rect 757 159 759 164
rect 769 159 771 164
rect 781 159 783 164
rect 793 160 795 164
rect 805 160 807 164
rect 817 160 819 164
rect 855 160 857 164
rect 894 160 896 164
rect 453 137 455 143
rect 208 55 210 66
rect 220 55 222 67
rect 254 55 256 66
rect 266 55 268 67
rect 288 56 290 60
rect -9 6 -7 12
rect 42 11 44 15
rect 54 12 56 15
rect 88 11 90 15
rect 100 12 102 15
rect 322 52 324 96
rect 334 72 336 96
rect 373 79 375 96
rect 419 79 421 96
rect 453 80 455 97
rect 704 90 706 95
rect 716 90 718 95
rect 728 90 730 95
rect 740 90 742 95
rect 752 90 754 95
rect 764 90 766 95
rect 776 90 778 95
rect 788 90 790 95
rect 826 90 828 95
rect 373 55 375 66
rect 385 55 387 67
rect 419 55 421 66
rect 431 55 433 67
rect 453 56 455 60
rect 157 6 159 12
rect 208 11 210 15
rect 220 12 222 15
rect 254 11 256 15
rect 266 12 268 15
rect 881 62 883 68
rect 322 6 324 12
rect 373 11 375 15
rect 385 12 387 15
rect 419 11 421 15
rect 431 12 433 15
rect 704 -14 706 50
rect 716 -14 718 50
rect -178 -75 -176 -71
rect -166 -75 -164 -71
rect -127 -75 -125 -71
rect -81 -75 -79 -71
rect -10 -75 -8 -71
rect 2 -75 4 -71
rect 41 -75 43 -71
rect 87 -75 89 -71
rect 156 -75 158 -71
rect 168 -75 170 -71
rect 207 -75 209 -71
rect 253 -75 255 -71
rect 321 -75 323 -71
rect 333 -75 335 -71
rect 372 -75 374 -71
rect 418 -75 420 -71
rect -47 -114 -45 -108
rect -178 -199 -176 -155
rect -166 -179 -164 -155
rect -127 -172 -125 -155
rect -81 -172 -79 -155
rect -47 -171 -45 -154
rect 121 -114 123 -108
rect -127 -196 -125 -185
rect -115 -196 -113 -184
rect -81 -196 -79 -185
rect -69 -196 -67 -184
rect -47 -195 -45 -191
rect -10 -199 -8 -155
rect 2 -179 4 -155
rect 41 -172 43 -155
rect 87 -172 89 -155
rect 121 -171 123 -154
rect 287 -114 289 -108
rect 41 -196 43 -185
rect 53 -196 55 -184
rect 87 -196 89 -185
rect 99 -196 101 -184
rect 121 -195 123 -191
rect -178 -245 -176 -239
rect -127 -240 -125 -236
rect -115 -239 -113 -236
rect -81 -240 -79 -236
rect -69 -239 -67 -236
rect 156 -199 158 -155
rect 168 -179 170 -155
rect 207 -172 209 -155
rect 253 -172 255 -155
rect 287 -171 289 -154
rect 704 -103 706 -18
rect 716 -103 718 -18
rect 728 -103 730 50
rect 740 -103 742 50
rect 752 -103 754 50
rect 764 -103 766 50
rect 776 -103 778 50
rect 788 -103 790 50
rect 826 -91 828 50
rect 881 5 883 22
rect 881 -19 883 -15
rect 452 -114 454 -108
rect 826 -115 828 -111
rect 704 -129 706 -123
rect 716 -126 718 -123
rect 728 -128 730 -123
rect 740 -127 742 -123
rect 752 -127 754 -123
rect 764 -128 766 -123
rect 776 -129 778 -123
rect 788 -128 790 -123
rect 207 -196 209 -185
rect 219 -196 221 -184
rect 253 -196 255 -185
rect 265 -196 267 -184
rect 287 -195 289 -191
rect -10 -245 -8 -239
rect 41 -240 43 -236
rect 53 -239 55 -236
rect 87 -240 89 -236
rect 99 -239 101 -236
rect 321 -199 323 -155
rect 333 -179 335 -155
rect 372 -172 374 -155
rect 418 -172 420 -155
rect 452 -171 454 -154
rect 372 -196 374 -185
rect 384 -196 386 -184
rect 418 -196 420 -185
rect 430 -196 432 -184
rect 452 -195 454 -191
rect 156 -245 158 -239
rect 207 -240 209 -236
rect 219 -239 221 -236
rect 253 -240 255 -236
rect 265 -239 267 -236
rect 321 -245 323 -239
rect 372 -240 374 -236
rect 384 -239 386 -236
rect 418 -240 420 -236
rect 430 -239 432 -236
rect 688 -268 690 -265
rect 700 -268 702 -265
rect 712 -268 714 -265
rect 724 -268 726 -265
rect 761 -268 763 -265
rect 793 -267 795 -261
rect 688 -350 690 -308
rect 700 -350 702 -308
rect 712 -350 714 -308
rect 724 -350 726 -308
rect 761 -350 763 -308
rect 688 -375 690 -370
rect 700 -375 702 -370
rect 712 -374 714 -370
rect 724 -374 726 -370
rect 761 -374 763 -370
rect 793 -373 795 -307
rect 793 -397 795 -393
<< polycontact >>
rect 702 796 707 802
rect 714 785 719 790
rect 733 777 738 782
rect 738 768 743 773
rect 750 758 755 764
rect 762 749 767 754
rect 774 741 779 746
rect 786 732 791 737
rect 798 723 803 728
rect 810 714 815 719
rect 822 705 827 710
rect 834 696 839 701
rect 846 687 851 692
rect 858 678 863 683
rect 870 669 875 674
rect 908 660 913 665
rect 947 651 952 656
rect 991 817 996 821
rect 693 360 697 364
rect 705 351 709 355
rect 723 343 727 347
rect 729 335 733 339
rect 741 325 745 329
rect 753 317 757 321
rect 765 309 769 313
rect 777 300 781 305
rect 789 290 793 295
rect 801 278 805 283
rect 813 268 817 273
rect 851 258 855 263
rect 890 249 894 254
rect 925 372 930 376
rect -183 67 -177 72
rect -51 83 -46 87
rect -163 75 -157 79
rect -128 75 -122 79
rect -82 75 -76 79
rect -127 66 -123 70
rect -115 67 -111 72
rect -81 66 -77 70
rect -69 67 -65 72
rect -15 67 -9 72
rect 117 83 122 87
rect 5 75 11 79
rect 40 75 46 79
rect 86 75 92 79
rect 41 66 45 70
rect 53 67 57 72
rect 87 66 91 70
rect 99 67 103 72
rect 151 67 157 72
rect 283 83 288 87
rect 171 75 177 79
rect 206 75 212 79
rect 252 75 258 79
rect 207 66 211 70
rect 219 67 223 72
rect 253 66 257 70
rect 265 67 269 72
rect 316 67 322 72
rect 448 83 453 87
rect 336 75 342 79
rect 371 75 377 79
rect 417 75 423 79
rect 372 66 376 70
rect 384 67 388 72
rect 418 66 422 70
rect 430 67 434 72
rect 700 -1 704 3
rect 712 -10 716 -6
rect 724 -18 728 -14
rect -184 -184 -178 -179
rect -52 -168 -47 -164
rect -164 -176 -158 -172
rect -129 -176 -123 -172
rect -83 -176 -77 -172
rect -128 -185 -124 -181
rect -116 -184 -112 -179
rect -82 -185 -78 -181
rect -70 -184 -66 -179
rect -16 -184 -10 -179
rect 116 -168 121 -164
rect 4 -176 10 -172
rect 39 -176 45 -172
rect 85 -176 91 -172
rect 40 -185 44 -181
rect 52 -184 56 -179
rect 86 -185 90 -181
rect 98 -184 102 -179
rect 150 -184 156 -179
rect 282 -168 287 -164
rect 736 -26 740 -22
rect 748 -34 752 -30
rect 760 -42 764 -38
rect 772 -52 776 -48
rect 784 -60 788 -56
rect 822 -68 826 -64
rect 876 9 881 13
rect 170 -176 176 -172
rect 205 -176 211 -172
rect 251 -176 257 -172
rect 206 -185 210 -181
rect 218 -184 222 -179
rect 252 -185 256 -181
rect 264 -184 268 -179
rect 315 -184 321 -179
rect 447 -168 452 -164
rect 335 -176 341 -172
rect 370 -176 376 -172
rect 416 -176 422 -172
rect 371 -185 375 -181
rect 383 -184 387 -179
rect 417 -185 421 -181
rect 429 -184 433 -179
rect 687 -265 691 -261
rect 699 -265 703 -261
rect 711 -265 715 -261
rect 723 -265 727 -261
rect 760 -265 764 -261
rect 788 -347 793 -343
<< metal1 >>
rect 525 942 994 946
rect 525 517 529 942
rect 702 929 706 942
rect 760 929 765 942
rect 844 929 849 942
rect 724 822 728 889
rect 736 833 741 889
rect 784 848 789 889
rect 796 871 801 889
rect 808 848 813 889
rect 819 868 824 889
rect 856 877 861 889
rect 867 887 872 889
rect 878 887 882 889
rect 909 877 912 889
rect 856 872 912 877
rect 916 868 920 889
rect 819 863 867 868
rect 872 863 920 868
rect 784 842 878 848
rect 736 829 795 833
rect 948 833 951 889
rect 802 829 951 833
rect 955 821 959 889
rect 991 870 994 942
rect 999 821 1003 830
rect 729 817 991 821
rect 999 817 1016 821
rect 724 808 728 813
rect 600 797 681 802
rect 595 796 681 797
rect 691 796 702 802
rect 662 785 714 790
rect 702 781 707 785
rect 702 777 733 781
rect 738 777 739 781
rect 702 776 739 777
rect 651 768 711 773
rect 717 768 738 773
rect 583 763 735 764
rect 588 758 735 763
rect 741 758 750 764
rect 574 749 698 754
rect 704 749 762 754
rect 641 741 747 746
rect 752 741 774 746
rect 717 732 786 737
rect 741 723 798 728
rect 752 714 810 719
rect 631 705 808 710
rect 813 705 822 710
rect 563 696 820 701
rect 826 696 834 701
rect 665 687 667 692
rect 673 687 846 692
rect 826 678 858 683
rect 704 669 870 674
rect 813 660 908 665
rect 680 651 681 656
rect 691 651 947 656
rect 736 639 794 645
rect 724 571 728 576
rect 736 571 741 639
rect 801 639 951 645
rect 784 626 878 631
rect 784 571 788 626
rect 795 571 800 583
rect 808 571 812 626
rect 819 596 867 603
rect 873 596 920 603
rect 819 571 823 596
rect 856 582 912 587
rect 856 571 860 582
rect 878 571 882 572
rect 908 571 912 582
rect 916 571 920 596
rect 947 571 951 639
rect 955 571 959 817
rect 999 813 1003 817
rect 702 541 706 551
rect 760 541 764 551
rect 844 541 848 551
rect 991 541 995 793
rect 701 536 995 541
rect 525 513 943 517
rect 525 190 529 513
rect 692 495 696 513
rect 750 495 754 513
rect 820 495 824 513
rect 714 376 718 455
rect 726 403 730 455
rect 774 426 778 455
rect 786 403 790 455
rect 798 426 802 455
rect 810 437 814 455
rect 851 437 854 455
rect 810 434 854 437
rect 858 427 862 455
rect 890 403 893 455
rect 726 399 893 403
rect 897 376 901 455
rect 925 425 928 513
rect 933 376 937 385
rect 719 372 925 376
rect 933 372 950 376
rect 719 371 901 372
rect 589 360 686 364
rect 692 360 693 364
rect 652 351 705 355
rect 692 347 696 351
rect 692 343 723 347
rect 727 343 729 347
rect 642 335 701 339
rect 706 335 729 339
rect 576 325 725 329
rect 731 325 741 329
rect 564 317 737 321
rect 742 317 753 321
rect 632 309 749 313
rect 755 309 765 313
rect 706 300 777 305
rect 731 290 789 295
rect 737 278 738 283
rect 743 278 801 283
rect 676 268 813 273
rect 755 258 851 263
rect 692 249 890 254
rect 726 233 893 237
rect -208 182 529 190
rect 714 184 718 227
rect 726 184 730 233
rect 774 184 777 204
rect 787 184 791 233
rect 799 184 802 205
rect 810 190 853 195
rect 810 184 813 190
rect 850 184 853 190
rect 858 184 861 205
rect 889 184 893 233
rect -208 -61 -197 182
rect -182 176 -178 182
rect -131 176 -127 182
rect -85 176 -81 182
rect -51 181 529 182
rect -51 137 -47 181
rect -14 176 -10 181
rect 37 176 41 181
rect 83 176 87 181
rect -162 86 -158 96
rect -174 82 -158 86
rect -123 87 -119 96
rect -136 83 -98 87
rect -77 87 -73 96
rect -43 88 -39 97
rect 117 137 121 181
rect 152 176 156 181
rect 203 176 207 181
rect 249 176 253 181
rect -90 83 -51 87
rect -43 84 -33 88
rect -27 84 -25 88
rect 6 86 10 96
rect -188 67 -183 72
rect -174 70 -170 82
rect -157 75 -151 79
rect -101 79 -98 83
rect -43 80 -39 84
rect -146 75 -128 79
rect -122 75 -104 79
rect -101 75 -82 79
rect -76 75 -65 79
rect -115 72 -111 75
rect -174 66 -127 70
rect -108 70 -104 75
rect -69 72 -65 75
rect -108 66 -81 70
rect -174 52 -170 66
rect -6 82 10 86
rect 45 87 49 96
rect 32 83 70 87
rect 91 87 95 96
rect 125 88 129 97
rect 283 137 287 181
rect 317 176 321 181
rect 368 176 372 181
rect 414 176 418 181
rect 78 83 117 87
rect 125 84 137 88
rect -20 67 -15 72
rect -6 70 -2 82
rect 11 75 17 79
rect 67 79 70 83
rect 125 80 129 84
rect 142 84 143 88
rect 172 86 176 96
rect 22 75 40 79
rect 46 75 64 79
rect 67 75 86 79
rect 92 75 103 79
rect 53 72 57 75
rect -6 66 41 70
rect 60 70 64 75
rect 99 72 103 75
rect 60 66 87 70
rect -182 6 -178 12
rect -111 6 -107 15
rect -65 6 -61 15
rect -51 6 -46 60
rect -6 52 -2 66
rect 160 82 176 86
rect 211 87 215 96
rect 198 83 236 87
rect 257 87 261 96
rect 291 88 295 97
rect 448 137 452 181
rect 244 83 283 87
rect 291 84 301 88
rect 146 67 151 72
rect 160 70 164 82
rect 177 75 183 79
rect 233 79 236 83
rect 291 80 295 84
rect 337 86 341 96
rect 188 75 206 79
rect 212 75 230 79
rect 233 75 252 79
rect 258 75 269 79
rect 219 72 223 75
rect 160 66 207 70
rect 226 70 230 75
rect 265 72 269 75
rect 226 66 253 70
rect -14 6 -10 12
rect 57 6 61 15
rect 103 6 107 15
rect 117 6 122 60
rect 160 52 164 66
rect 325 82 341 86
rect 376 87 380 96
rect 363 83 401 87
rect 422 87 426 96
rect 456 88 460 97
rect 525 110 529 181
rect 897 184 901 371
rect 933 368 937 372
rect 692 143 696 164
rect 750 143 754 164
rect 820 143 824 164
rect 925 143 929 348
rect 991 143 995 536
rect 692 138 995 143
rect 525 106 879 110
rect 409 83 448 87
rect 456 84 470 88
rect 311 67 316 72
rect 325 70 329 82
rect 342 75 348 79
rect 398 79 401 83
rect 456 80 460 84
rect 353 75 371 79
rect 377 75 395 79
rect 398 75 417 79
rect 423 75 434 79
rect 384 72 388 75
rect 325 66 372 70
rect 391 70 395 75
rect 430 72 434 75
rect 391 66 418 70
rect 152 6 156 12
rect 223 6 227 15
rect 269 6 273 15
rect 283 6 288 60
rect 325 52 329 66
rect 317 6 321 12
rect 388 6 392 15
rect 434 6 438 15
rect 448 6 453 60
rect -186 1 502 6
rect -208 -69 451 -61
rect -183 -75 -179 -69
rect -132 -75 -128 -69
rect -86 -75 -82 -69
rect -52 -70 451 -69
rect -52 -114 -48 -70
rect -15 -75 -11 -70
rect 36 -75 40 -70
rect 82 -75 86 -70
rect -163 -165 -159 -155
rect -175 -169 -159 -165
rect -124 -164 -120 -155
rect -137 -168 -99 -164
rect -78 -164 -74 -155
rect -44 -163 -40 -154
rect 116 -114 120 -70
rect 151 -75 155 -70
rect 202 -75 206 -70
rect 248 -75 252 -70
rect -91 -168 -52 -164
rect -44 -167 -34 -163
rect -28 -167 -26 -163
rect 5 -165 9 -155
rect -189 -184 -184 -179
rect -175 -181 -171 -169
rect -158 -176 -152 -172
rect -102 -172 -99 -168
rect -44 -171 -40 -167
rect -147 -176 -129 -172
rect -123 -176 -105 -172
rect -102 -176 -83 -172
rect -77 -176 -66 -172
rect -116 -179 -112 -176
rect -175 -185 -128 -181
rect -109 -181 -105 -176
rect -70 -179 -66 -176
rect -109 -185 -82 -181
rect -175 -199 -171 -185
rect -7 -169 9 -165
rect 44 -164 48 -155
rect 31 -168 69 -164
rect 90 -164 94 -155
rect 124 -163 128 -154
rect 282 -114 286 -70
rect 316 -75 320 -70
rect 367 -75 371 -70
rect 413 -75 417 -70
rect 77 -168 116 -164
rect 124 -167 136 -163
rect -21 -184 -16 -179
rect -7 -181 -3 -169
rect 10 -176 16 -172
rect 66 -172 69 -168
rect 124 -171 128 -167
rect 141 -167 142 -163
rect 171 -165 175 -155
rect 21 -176 39 -172
rect 45 -176 63 -172
rect 66 -176 85 -172
rect 91 -176 102 -172
rect 52 -179 56 -176
rect -7 -185 40 -181
rect 59 -181 63 -176
rect 98 -179 102 -176
rect 59 -185 86 -181
rect -183 -245 -179 -239
rect -112 -245 -108 -236
rect -66 -245 -62 -236
rect -52 -245 -47 -191
rect -7 -199 -3 -185
rect 159 -169 175 -165
rect 210 -164 214 -155
rect 197 -168 235 -164
rect 256 -164 260 -155
rect 290 -163 294 -154
rect 447 -114 451 -70
rect 243 -168 282 -164
rect 290 -167 300 -163
rect 145 -184 150 -179
rect 159 -181 163 -169
rect 176 -176 182 -172
rect 232 -172 235 -168
rect 290 -171 294 -167
rect 336 -165 340 -155
rect 187 -176 205 -172
rect 211 -176 229 -172
rect 232 -176 251 -172
rect 257 -176 268 -172
rect 218 -179 222 -176
rect 159 -185 206 -181
rect 225 -181 229 -176
rect 264 -179 268 -176
rect 225 -185 252 -181
rect -15 -245 -11 -239
rect 56 -245 60 -236
rect 102 -245 106 -236
rect 116 -245 121 -191
rect 159 -199 163 -185
rect 324 -169 340 -165
rect 375 -164 379 -155
rect 362 -168 400 -164
rect 421 -164 425 -155
rect 455 -163 459 -154
rect 408 -168 447 -164
rect 455 -167 469 -163
rect 310 -184 315 -179
rect 324 -181 328 -169
rect 341 -176 347 -172
rect 397 -172 400 -168
rect 455 -171 459 -167
rect 352 -176 370 -172
rect 376 -176 394 -172
rect 397 -176 416 -172
rect 422 -176 433 -172
rect 383 -179 387 -176
rect 324 -185 371 -181
rect 390 -181 394 -176
rect 429 -179 433 -176
rect 390 -185 417 -181
rect 151 -245 155 -239
rect 222 -245 226 -236
rect 268 -245 272 -236
rect 282 -245 287 -191
rect 324 -199 328 -185
rect 316 -245 320 -239
rect 387 -245 391 -236
rect 433 -245 437 -236
rect 447 -245 452 -191
rect 497 -245 502 1
rect 525 -211 529 106
rect 558 99 564 100
rect 558 58 564 94
rect 570 99 576 100
rect 570 68 576 94
rect 583 78 589 93
rect 699 90 703 106
rect 757 90 761 106
rect 769 98 825 101
rect 769 90 773 98
rect 821 90 825 98
rect 721 14 724 50
rect 733 21 736 50
rect 782 21 785 50
rect 791 39 794 50
rect 829 21 833 50
rect 876 62 879 106
rect 733 18 833 21
rect 725 10 791 13
rect 884 13 888 22
rect 796 10 876 13
rect 884 9 904 13
rect 721 7 724 9
rect 884 5 888 9
rect 577 -1 680 3
rect 686 -1 700 3
rect 641 -10 712 -6
rect 699 -14 702 -10
rect 699 -18 724 -14
rect 632 -26 708 -22
rect 713 -26 736 -22
rect 564 -34 691 -30
rect 696 -34 748 -30
rect 675 -42 760 -38
rect 696 -52 772 -48
rect 686 -60 784 -56
rect 713 -68 822 -64
rect 733 -78 833 -75
rect 721 -103 724 -79
rect 733 -103 736 -78
rect 781 -103 784 -78
rect 791 -103 794 -86
rect 830 -91 833 -78
rect 699 -140 703 -123
rect 770 -132 773 -123
rect 821 -132 824 -111
rect 770 -135 824 -132
rect 876 -140 880 -15
rect 925 -140 929 138
rect 699 -143 929 -140
rect 699 -145 880 -143
rect 544 -166 607 -163
rect 544 -167 617 -166
rect 547 -179 610 -174
rect 616 -179 618 -174
rect 547 -189 608 -184
rect 617 -189 618 -184
rect 626 -194 631 -159
rect 636 -184 641 -159
rect 646 -173 652 -158
rect 547 -199 610 -194
rect 525 -216 786 -211
rect 564 -226 727 -222
rect 632 -238 691 -234
rect 687 -241 691 -238
rect -187 -250 502 -245
rect 447 -400 452 -250
rect 687 -261 691 -246
rect 699 -261 703 -255
rect 711 -261 715 -237
rect 723 -250 727 -226
rect 723 -261 727 -255
rect 760 -261 764 -246
rect 782 -257 786 -216
rect 782 -261 806 -257
rect 788 -267 792 -261
rect 731 -303 736 -299
rect 683 -324 687 -308
rect 683 -350 687 -329
rect 705 -334 709 -308
rect 717 -317 720 -308
rect 757 -317 760 -308
rect 717 -321 760 -317
rect 764 -325 768 -308
rect 764 -343 768 -330
rect 788 -333 792 -307
rect 796 -343 800 -307
rect 764 -347 788 -343
rect 796 -347 816 -343
rect 764 -350 768 -347
rect 731 -363 735 -359
rect 683 -390 687 -370
rect 693 -376 697 -370
rect 705 -400 709 -370
rect 717 -380 721 -370
rect 756 -380 760 -370
rect 717 -384 760 -380
rect 764 -389 768 -370
rect 796 -373 800 -347
rect 788 -400 793 -393
rect 876 -400 880 -145
rect 447 -404 880 -400
rect 868 -405 879 -404
<< m2contact >>
rect 795 865 802 871
rect 867 881 872 887
rect 878 881 884 887
rect 867 862 872 868
rect 878 840 884 849
rect 795 828 802 834
rect 723 813 729 822
rect 595 797 600 802
rect 681 794 691 802
rect 657 785 662 790
rect 646 768 651 773
rect 711 768 717 773
rect 583 758 588 763
rect 735 758 741 764
rect 569 749 574 754
rect 698 749 704 754
rect 636 741 641 746
rect 747 741 752 746
rect 711 732 717 737
rect 735 723 741 729
rect 747 714 752 719
rect 626 705 631 710
rect 808 705 813 710
rect 558 696 563 701
rect 820 696 826 701
rect 667 687 673 692
rect 820 678 826 683
rect 698 669 704 674
rect 808 660 813 665
rect 681 650 691 658
rect 723 576 729 585
rect 794 638 801 646
rect 794 583 802 591
rect 878 625 883 632
rect 867 596 873 603
rect 867 571 873 578
rect 878 572 883 577
rect 773 421 779 426
rect 797 421 803 426
rect 858 422 864 427
rect 713 370 719 376
rect 583 360 589 365
rect 686 359 692 365
rect 646 351 652 356
rect 636 335 642 340
rect 701 334 706 340
rect 570 324 576 329
rect 725 324 731 330
rect 558 316 564 321
rect 737 317 742 322
rect 626 309 632 314
rect 749 308 755 314
rect 701 299 706 306
rect 725 289 731 296
rect 738 278 743 283
rect 667 268 676 273
rect 749 257 755 263
rect 686 248 692 254
rect 713 227 718 232
rect 773 204 778 209
rect 799 205 804 210
rect 858 205 863 210
rect -141 83 -136 88
rect -95 83 -90 88
rect -33 84 -27 90
rect -151 75 -146 80
rect 27 83 32 88
rect 73 83 78 88
rect 17 75 22 80
rect 137 83 142 88
rect -132 55 -127 60
rect -86 55 -81 60
rect 193 83 198 88
rect 239 83 244 88
rect 183 75 188 80
rect 301 83 306 89
rect 36 55 41 60
rect 82 55 87 60
rect 358 83 363 88
rect 404 83 409 88
rect 348 75 353 80
rect 470 83 476 89
rect 202 55 207 60
rect 248 55 253 60
rect 367 55 372 60
rect 413 55 418 60
rect -142 -168 -137 -163
rect -96 -168 -91 -163
rect -34 -167 -28 -161
rect -152 -176 -147 -171
rect 26 -168 31 -163
rect 72 -168 77 -163
rect 16 -176 21 -171
rect 136 -168 141 -163
rect -133 -196 -128 -191
rect -87 -196 -82 -191
rect 192 -168 197 -163
rect 238 -168 243 -163
rect 182 -176 187 -171
rect 300 -168 305 -162
rect 35 -196 40 -191
rect 81 -196 86 -191
rect 357 -168 362 -163
rect 403 -168 408 -163
rect 347 -176 352 -171
rect 469 -168 475 -162
rect 201 -196 206 -191
rect 247 -196 252 -191
rect 366 -196 371 -191
rect 412 -196 417 -191
rect 557 94 564 99
rect 570 94 577 99
rect 583 93 590 98
rect 583 72 590 78
rect 570 62 577 68
rect 558 52 565 58
rect 791 33 796 39
rect 720 9 725 14
rect 791 9 796 14
rect 569 -2 577 3
rect 680 -1 686 4
rect 635 -11 641 -5
rect 626 -26 632 -20
rect 708 -26 713 -21
rect 558 -35 564 -29
rect 691 -34 696 -29
rect 667 -42 675 -37
rect 691 -52 696 -47
rect 680 -60 686 -55
rect 708 -68 713 -63
rect 720 -79 725 -74
rect 791 -86 796 -81
rect 625 -159 631 -154
rect 635 -159 642 -154
rect 646 -158 652 -152
rect 538 -168 544 -161
rect 607 -166 617 -161
rect 538 -179 547 -174
rect 610 -179 616 -172
rect 538 -189 547 -184
rect 608 -189 617 -184
rect 645 -180 653 -173
rect 634 -190 641 -184
rect 538 -199 547 -194
rect 610 -199 619 -194
rect 625 -200 631 -194
rect 557 -227 564 -222
rect 624 -239 632 -234
rect 710 -237 716 -232
rect 686 -246 691 -241
rect 699 -255 704 -250
rect 759 -246 764 -241
rect 722 -255 727 -250
rect 736 -303 742 -298
rect 681 -329 687 -324
rect 704 -339 709 -334
rect 764 -330 770 -325
rect 787 -339 792 -333
rect 735 -364 740 -357
rect 683 -396 688 -390
rect 763 -396 770 -389
<< metal2 >>
rect 867 868 872 881
rect 796 834 801 865
rect 878 849 882 881
rect 558 701 564 812
rect 570 754 576 812
rect 574 749 576 754
rect 563 696 564 701
rect 558 321 564 696
rect -228 195 353 199
rect -228 -51 -223 195
rect -151 80 -146 195
rect -151 74 -146 75
rect -141 60 -136 83
rect -95 60 -90 83
rect -141 55 -132 60
rect -95 55 -86 60
rect -32 -23 -28 84
rect 17 80 22 195
rect 27 60 32 83
rect 73 60 78 83
rect 27 55 36 60
rect 73 55 82 60
rect 137 -13 141 83
rect 183 80 188 195
rect 193 60 198 83
rect 239 60 244 83
rect 193 55 202 60
rect 239 55 248 60
rect 301 -4 305 83
rect 348 80 353 195
rect 558 99 564 316
rect 570 329 576 749
rect 570 99 576 324
rect 583 763 589 812
rect 588 758 589 763
rect 583 365 589 758
rect 583 98 589 360
rect 595 802 600 812
rect 358 60 363 83
rect 595 88 600 797
rect 476 84 600 88
rect 404 60 409 83
rect 473 72 583 77
rect 358 55 367 60
rect 404 55 413 60
rect 473 -4 478 72
rect 301 -8 478 -4
rect 487 62 570 67
rect 487 -13 491 62
rect 137 -17 491 -13
rect 497 52 558 57
rect 497 -23 501 52
rect -32 -28 501 -23
rect 558 -29 564 52
rect 570 3 576 62
rect -228 -56 351 -51
rect -152 -171 -148 -56
rect -142 -191 -137 -168
rect -96 -191 -91 -168
rect -142 -196 -133 -191
rect -96 -196 -87 -191
rect -33 -274 -29 -167
rect 16 -171 20 -56
rect 26 -191 31 -168
rect 72 -191 77 -168
rect 26 -196 35 -191
rect 72 -196 81 -191
rect 136 -264 140 -168
rect 182 -171 186 -56
rect 346 -57 351 -56
rect 192 -191 197 -168
rect 238 -191 243 -168
rect 192 -196 201 -191
rect 238 -196 247 -191
rect 300 -255 304 -168
rect 347 -171 351 -57
rect 357 -191 362 -168
rect 475 -167 538 -163
rect 403 -191 408 -168
rect 472 -179 538 -174
rect 357 -196 366 -191
rect 403 -196 412 -191
rect 472 -255 477 -179
rect 300 -259 477 -255
rect 486 -189 538 -184
rect 486 -264 490 -189
rect 136 -268 490 -264
rect 496 -199 538 -194
rect 496 -274 500 -199
rect 558 -222 564 -35
rect 558 -249 564 -227
rect 570 -249 576 -2
rect 583 -249 589 72
rect 595 -249 600 84
rect 626 710 631 812
rect 626 314 631 705
rect 636 746 641 812
rect 636 340 641 741
rect 646 773 652 812
rect 651 768 652 773
rect 646 356 652 768
rect 626 -20 631 309
rect 636 -5 641 335
rect 626 -154 631 -26
rect 636 -154 641 -11
rect 646 -152 652 351
rect 657 790 662 812
rect 657 -163 662 785
rect 617 -166 662 -163
rect 607 -167 662 -166
rect 608 -179 610 -174
rect 616 -179 645 -174
rect 617 -189 634 -184
rect 608 -199 610 -194
rect 619 -199 625 -194
rect 626 -234 631 -200
rect 626 -249 631 -239
rect 636 -249 641 -190
rect 646 -249 652 -180
rect 657 -249 662 -167
rect 667 273 673 687
rect 682 658 690 794
rect 698 674 704 749
rect 711 737 717 768
rect 724 585 728 813
rect 735 729 741 758
rect 747 719 752 741
rect 808 665 812 705
rect 820 683 825 696
rect 795 591 800 638
rect 868 578 872 596
rect 724 571 728 576
rect 878 577 882 625
rect 878 571 882 572
rect 779 422 797 426
rect 803 422 858 426
rect 714 376 718 377
rect 667 -37 675 268
rect 686 254 692 359
rect 701 306 705 334
rect 714 232 718 370
rect 726 296 730 324
rect 742 317 743 321
rect 737 283 743 317
rect 737 278 738 283
rect 750 263 754 308
rect 778 205 799 209
rect 804 205 858 209
rect 791 14 794 33
rect 667 -202 675 -42
rect 681 -55 686 -1
rect 721 -14 724 9
rect 692 -47 696 -34
rect 709 -63 713 -26
rect 721 -74 724 -18
rect 791 -81 794 9
rect 791 -91 794 -86
rect 667 -206 715 -202
rect 711 -232 715 -206
rect 691 -246 759 -242
rect 704 -255 722 -251
rect -33 -279 500 -274
rect 736 -326 741 -303
rect 687 -329 764 -326
rect 709 -339 787 -334
rect 735 -391 739 -364
rect 688 -395 763 -391
<< labels >>
rlabel metal1 -154 77 -154 77 1 clk
rlabel metal1 -174 2 -174 2 1 gnd
rlabel metal1 -81 187 -81 187 5 vdd
rlabel metal1 -127 187 -127 187 5 vdd
rlabel metal1 -170 188 -170 188 5 vdd
rlabel metal1 -187 68 -185 71 3 a0_in
rlabel metal1 -36 85 -33 87 1 a0
rlabel metal1 14 77 14 77 1 clk
rlabel metal1 -6 2 -6 2 1 gnd
rlabel metal1 87 187 87 187 5 vdd
rlabel metal1 41 187 41 187 5 vdd
rlabel metal1 -2 188 -2 188 5 vdd
rlabel metal1 -20 67 -14 72 1 a1_in
rlabel metal1 132 84 136 88 1 a1
rlabel metal1 180 77 180 77 1 clk
rlabel metal1 160 2 160 2 1 gnd
rlabel metal1 253 187 253 187 5 vdd
rlabel metal1 207 187 207 187 5 vdd
rlabel metal1 164 188 164 188 5 vdd
rlabel space 146 67 152 73 1 a2_in
rlabel space 298 83 303 89 1 a2
rlabel metal1 345 77 345 77 1 clk
rlabel metal1 325 2 325 2 1 gnd
rlabel metal1 418 187 418 187 5 vdd
rlabel metal1 372 187 372 187 5 vdd
rlabel metal1 329 188 329 188 5 vdd
rlabel metal1 311 67 316 72 1 a3_in
rlabel metal1 463 84 467 88 1 a3
rlabel metal2 503 84 508 88 1 a3
rlabel metal2 504 73 508 77 1 a2
rlabel space 504 61 509 67 1 a1
rlabel metal1 -155 -174 -155 -174 1 clk
rlabel metal1 -175 -249 -175 -249 1 gnd
rlabel metal1 -82 -64 -82 -64 5 vdd
rlabel metal1 -128 -64 -128 -64 5 vdd
rlabel metal1 -171 -63 -171 -63 5 vdd
rlabel metal1 13 -174 13 -174 1 clk
rlabel metal1 -7 -249 -7 -249 1 gnd
rlabel metal1 86 -64 86 -64 5 vdd
rlabel metal1 40 -64 40 -64 5 vdd
rlabel metal1 -3 -63 -3 -63 5 vdd
rlabel metal1 179 -174 179 -174 1 clk
rlabel metal1 159 -249 159 -249 1 gnd
rlabel metal1 252 -64 252 -64 5 vdd
rlabel metal1 206 -64 206 -64 5 vdd
rlabel metal1 163 -63 163 -63 5 vdd
rlabel metal1 344 -174 344 -174 1 clk
rlabel metal1 324 -249 324 -249 1 gnd
rlabel metal1 417 -64 417 -64 5 vdd
rlabel metal1 371 -64 371 -64 5 vdd
rlabel metal1 328 -63 328 -63 5 vdd
rlabel metal1 -189 -184 -182 -179 3 b0_in
rlabel space -38 -168 -34 -163 1 b0
rlabel metal1 -21 -184 -15 -179 1 b1_in
rlabel space 131 -168 135 -162 1 b1
rlabel metal1 145 -184 150 -179 1 b2_in
rlabel metal1 296 -167 299 -163 1 b2
rlabel metal1 310 -184 315 -179 1 b3_in
rlabel metal1 462 -167 466 -163 1 b3
rlabel metal2 498 -167 503 -163 1 b3
rlabel metal2 498 -178 503 -174 1 b2
rlabel metal2 498 -189 503 -185 1 b1
rlabel metal2 501 -199 506 -195 1 b0
rlabel metal1 668 -26 674 -22 1 b0
rlabel m2contact 669 -42 674 -38 1 cin
rlabel metal1 668 -34 673 -30 1 a0
rlabel metal1 668 -1 672 3 1 a1
rlabel metal1 930 516 930 516 5 vdd
rlabel metal1 681 360 686 364 1 a2
rlabel metal1 682 351 687 355 1 b2
rlabel metal1 683 335 687 339 1 b1
rlabel metal1 683 325 687 329 1 a1
rlabel metal1 684 317 688 321 1 a0
rlabel metal1 685 309 689 313 1 b0
rlabel metal1 685 268 690 273 1 cin
rlabel metal1 942 372 949 376 7 c3
rlabel metal1 930 141 930 141 1 gnd
rlabel metal1 670 797 675 802 1 a3
rlabel metal1 670 768 676 773 1 b2
rlabel metal1 670 759 676 764 1 a2
rlabel metal1 670 741 676 746 1 b1
rlabel metal1 666 785 671 790 1 b3
rlabel metal1 666 749 671 754 1 a1
rlabel metal1 675 706 680 710 1 b0
rlabel metal1 676 696 681 700 1 a0
rlabel metal1 675 687 681 692 1 cin
rlabel metal1 686 -10 692 -6 3 b1
rlabel metal1 726 -144 732 -142 1 gnd
rlabel metal1 728 107 732 109 5 vdd
rlabel metal1 892 9 897 13 1 c2
rlabel metal1 869 107 878 110 5 vdd
rlabel metal1 858 -145 866 -140 1 gnd
rlabel metal1 1007 817 1012 821 1 cout
rlabel metal1 956 942 963 945 5 vdd
rlabel space 521 52 526 58 1 a0
rlabel metal1 689 -259 689 -259 1 b0
rlabel metal1 702 -259 702 -259 1 a0
rlabel metal1 713 -259 713 -259 1 cin
rlabel metal1 725 -259 725 -259 1 a0
rlabel metal1 763 -259 763 -259 1 b0
rlabel metal1 793 -259 793 -259 5 vdd
rlabel metal1 684 -331 684 -331 1 n010
rlabel metal2 741 -328 741 -328 1 n010
rlabel metal1 793 -402 793 -402 1 gnd
rlabel metal2 738 -393 738 -393 1 n010
rlabel metal1 777 -345 777 -345 1 n010
rlabel metal1 809 -345 809 -345 1 c1
rlabel metal1 707 -381 707 -381 1 gnd
<< end >>
