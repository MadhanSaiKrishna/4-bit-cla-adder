magic
tech scmos
timestamp 1733201153
<< nwell >>
rect 349 81 457 133
rect 471 81 495 133
rect 526 53 550 105
<< ntransistor >>
rect 537 22 539 42
rect 360 -86 362 -66
rect 372 -86 374 -66
rect 384 -86 386 -66
rect 396 -86 398 -66
rect 408 -86 410 -66
rect 420 -86 422 -66
rect 432 -86 434 -66
rect 444 -86 446 -66
rect 482 -74 484 -54
<< ptransistor >>
rect 360 87 362 127
rect 372 87 374 127
rect 384 87 386 127
rect 396 87 398 127
rect 408 87 410 127
rect 420 87 422 127
rect 432 87 434 127
rect 444 87 446 127
rect 482 87 484 127
rect 537 59 539 99
<< ndiffusion >>
rect 536 22 537 42
rect 539 22 540 42
rect 359 -86 360 -66
rect 362 -86 363 -66
rect 371 -86 372 -66
rect 374 -86 375 -66
rect 383 -86 384 -66
rect 386 -86 387 -66
rect 395 -86 396 -66
rect 398 -86 399 -66
rect 407 -86 408 -66
rect 410 -86 411 -66
rect 419 -86 420 -66
rect 422 -86 423 -66
rect 431 -86 432 -66
rect 434 -86 435 -66
rect 443 -86 444 -66
rect 446 -86 447 -66
rect 481 -74 482 -54
rect 484 -74 485 -54
<< pdiffusion >>
rect 359 87 360 127
rect 362 87 363 127
rect 371 87 372 127
rect 374 87 375 127
rect 383 87 384 127
rect 386 87 387 127
rect 395 87 396 127
rect 398 87 399 127
rect 407 87 408 127
rect 410 87 411 127
rect 419 87 420 127
rect 422 87 423 127
rect 431 87 432 127
rect 434 87 435 127
rect 443 87 444 127
rect 446 87 447 127
rect 481 87 482 127
rect 484 87 485 127
rect 536 59 537 99
rect 539 59 540 99
<< ndcontact >>
rect 532 22 536 42
rect 540 22 544 42
rect 355 -86 359 -66
rect 363 -86 371 -66
rect 375 -86 383 -66
rect 387 -86 395 -66
rect 399 -86 407 -66
rect 411 -86 419 -66
rect 423 -86 431 -66
rect 435 -86 443 -66
rect 447 -86 451 -66
rect 477 -74 481 -54
rect 485 -74 489 -54
<< pdcontact >>
rect 355 87 359 127
rect 363 87 371 127
rect 375 87 383 127
rect 387 87 395 127
rect 399 87 407 127
rect 411 87 419 127
rect 423 87 431 127
rect 435 87 443 127
rect 447 87 451 127
rect 477 87 481 127
rect 485 87 489 127
rect 532 59 536 99
rect 540 59 544 99
<< polysilicon >>
rect 360 127 362 132
rect 372 127 374 132
rect 384 127 386 132
rect 396 127 398 132
rect 408 127 410 132
rect 420 127 422 132
rect 432 127 434 132
rect 444 127 446 132
rect 482 127 484 132
rect 537 99 539 105
rect 360 23 362 87
rect 372 23 374 87
rect 360 -66 362 19
rect 372 -66 374 19
rect 384 -66 386 87
rect 396 -66 398 87
rect 408 -66 410 87
rect 420 -66 422 87
rect 432 -66 434 87
rect 444 -66 446 87
rect 482 -54 484 87
rect 537 42 539 59
rect 537 18 539 22
rect 482 -78 484 -74
rect 360 -92 362 -86
rect 372 -89 374 -86
rect 384 -91 386 -86
rect 396 -90 398 -86
rect 408 -90 410 -86
rect 420 -91 422 -86
rect 432 -92 434 -86
rect 444 -91 446 -86
<< polycontact >>
rect 356 36 360 40
rect 368 27 372 31
rect 380 19 384 23
rect 392 11 396 15
rect 404 3 408 7
rect 416 -5 420 -1
rect 428 -15 432 -11
rect 440 -23 444 -19
rect 478 -31 482 -27
rect 532 46 537 50
<< metal1 >>
rect 355 143 535 147
rect 355 127 359 143
rect 413 127 417 143
rect 425 135 481 138
rect 425 127 429 135
rect 477 127 481 135
rect 377 51 380 87
rect 389 58 392 87
rect 438 58 441 87
rect 447 76 450 87
rect 485 58 489 87
rect 532 99 535 143
rect 389 55 489 58
rect 381 47 447 50
rect 540 50 544 59
rect 452 47 532 50
rect 540 46 560 50
rect 377 44 380 46
rect 540 42 544 46
rect 326 36 336 40
rect 342 36 356 40
rect 326 27 368 31
rect 355 23 358 27
rect 355 19 380 23
rect 327 11 364 15
rect 369 11 392 15
rect 327 3 347 7
rect 352 3 404 7
rect 327 -5 416 -1
rect 352 -15 428 -11
rect 342 -23 440 -19
rect 369 -31 478 -27
rect 389 -41 489 -38
rect 377 -66 380 -42
rect 389 -66 392 -41
rect 437 -66 440 -41
rect 447 -66 450 -49
rect 486 -54 489 -41
rect 355 -103 359 -86
rect 426 -95 429 -86
rect 477 -95 480 -74
rect 426 -98 480 -95
rect 532 -103 536 22
rect 355 -108 536 -103
<< m2contact >>
rect 447 70 452 76
rect 376 46 381 51
rect 447 46 452 51
rect 336 36 342 41
rect 364 11 369 16
rect 347 3 352 8
rect 347 -15 352 -10
rect 336 -23 342 -18
rect 364 -31 369 -26
rect 376 -42 381 -37
rect 447 -49 452 -44
<< metal2 >>
rect 447 51 450 70
rect 337 -18 342 36
rect 377 23 380 46
rect 348 -10 352 3
rect 365 -26 369 11
rect 377 -37 380 19
rect 447 -44 450 46
rect 447 -54 450 -49
<< labels >>
rlabel metal1 328 27 334 31 3 b1
rlabel metal1 330 11 336 15 1 b0
rlabel metal1 331 -5 336 -1 1 cin
rlabel metal1 330 3 335 7 1 a0
rlabel metal1 382 -107 388 -105 1 gnd
rlabel metal1 384 144 388 146 5 vdd
rlabel metal1 330 36 334 40 1 a1
rlabel metal1 548 46 553 50 1 c2
rlabel metal1 525 144 534 147 5 vdd
rlabel metal1 514 -108 522 -103 1 gnd
<< end >>
