magic
tech scmos
timestamp 1733165166
<< nwell >>
rect 349 160 458 213
rect 471 160 496 213
rect 540 139 564 191
<< ntransistor >>
rect 551 108 553 128
rect 360 87 362 107
rect 372 87 374 107
rect 384 87 386 107
rect 396 87 398 107
rect 408 87 410 107
rect 420 87 422 107
rect 432 87 434 107
rect 444 87 446 107
rect 482 87 484 107
<< ptransistor >>
rect 360 166 362 206
rect 372 166 374 206
rect 384 166 386 206
rect 396 166 398 206
rect 408 166 410 206
rect 420 166 422 206
rect 432 166 434 206
rect 444 166 446 206
rect 482 166 484 206
rect 551 145 553 185
<< ndiffusion >>
rect 550 108 551 128
rect 553 108 554 128
rect 359 87 360 107
rect 362 87 363 107
rect 371 87 372 107
rect 374 87 375 107
rect 383 87 384 107
rect 386 87 387 107
rect 395 87 396 107
rect 398 87 399 107
rect 407 87 408 107
rect 410 87 411 107
rect 419 87 420 107
rect 422 87 423 107
rect 431 87 432 107
rect 434 87 435 107
rect 443 87 444 107
rect 446 87 447 107
rect 481 87 482 107
rect 484 87 485 107
<< pdiffusion >>
rect 359 166 360 206
rect 362 166 363 206
rect 371 166 372 206
rect 374 166 375 206
rect 383 166 384 206
rect 386 166 387 206
rect 395 166 396 206
rect 398 166 399 206
rect 407 166 408 206
rect 410 166 411 206
rect 419 166 420 206
rect 422 166 423 206
rect 431 166 432 206
rect 434 166 435 206
rect 443 166 444 206
rect 446 166 447 206
rect 481 166 482 206
rect 484 166 485 206
rect 550 145 551 185
rect 553 145 554 185
<< ndcontact >>
rect 546 108 550 128
rect 554 108 558 128
rect 355 87 359 107
rect 363 87 371 107
rect 375 87 383 107
rect 387 87 395 107
rect 399 87 407 107
rect 411 87 419 107
rect 423 87 431 107
rect 435 87 443 107
rect 447 87 451 107
rect 477 87 481 107
rect 485 87 489 107
<< pdcontact >>
rect 355 166 359 206
rect 363 166 371 206
rect 375 166 383 206
rect 387 166 395 206
rect 399 166 407 206
rect 411 166 419 206
rect 423 166 431 206
rect 435 166 443 206
rect 447 166 451 206
rect 477 166 481 206
rect 485 166 489 206
rect 546 145 550 185
rect 554 145 558 185
<< polysilicon >>
rect 360 206 362 209
rect 372 206 374 209
rect 384 206 386 209
rect 396 206 398 209
rect 408 206 410 209
rect 420 206 422 209
rect 432 206 434 209
rect 444 206 446 209
rect 482 206 484 209
rect 551 185 553 191
rect 360 107 362 166
rect 372 107 374 166
rect 384 107 386 166
rect 396 107 398 166
rect 408 107 410 166
rect 420 107 422 166
rect 432 107 434 166
rect 444 107 446 166
rect 482 107 484 166
rect 551 128 553 145
rect 551 104 553 108
rect 360 83 362 87
rect 372 83 374 87
rect 384 82 386 87
rect 396 82 398 87
rect 408 82 410 87
rect 420 83 422 87
rect 432 83 434 87
rect 444 83 446 87
rect 482 83 484 87
<< polycontact >>
rect 359 209 363 213
rect 371 209 375 213
rect 383 209 387 213
rect 395 209 399 213
rect 407 209 411 213
rect 419 209 423 213
rect 431 209 435 213
rect 443 209 447 213
rect 481 209 485 213
rect 546 132 551 136
<< metal1 >>
rect 359 213 363 223
rect 371 213 375 223
rect 383 213 387 223
rect 395 213 399 219
rect 407 213 411 223
rect 419 213 423 231
rect 431 213 435 231
rect 443 213 447 232
rect 481 213 485 219
rect 401 155 405 166
rect 413 158 417 166
rect 425 158 428 166
rect 478 158 481 166
rect 540 191 564 195
rect 485 158 489 166
rect 546 185 550 191
rect 554 136 558 145
rect 532 132 546 136
rect 554 132 574 136
rect 554 128 558 132
rect 485 107 489 110
rect 355 82 359 87
rect 377 80 381 87
rect 391 80 395 87
rect 401 81 405 87
rect 425 80 429 87
rect 477 80 481 87
rect 546 104 551 108
rect 540 100 564 104
rect 485 80 489 87
<< labels >>
rlabel metal1 397 215 397 215 1 b0
rlabel metal1 410 215 410 215 1 a0
rlabel metal1 421 215 421 215 1 cin
rlabel metal1 433 215 433 215 1 a0
rlabel metal1 445 218 445 218 1 a1
rlabel metal1 484 215 484 215 1 b0
rlabel metal1 373 218 373 218 1 b1
rlabel metal1 385 219 385 219 1 b1
rlabel metal1 359 217 362 220 1 a1
rlabel metal1 551 193 551 193 5 vdd
rlabel metal1 551 102 551 102 1 gnd
<< end >>
